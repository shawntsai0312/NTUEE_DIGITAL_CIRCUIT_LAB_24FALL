module Top (
	input i_rst_n,
	input i_clk,
	input i_key_0, // reset
	input i_key_1, // start
	input i_key_2, // stop
	input [3:0] i_speed, // design how user can decide mode on your own
	
	// AudDSP and SRAM
	output [19:0] o_SRAM_ADDR,
	inout  [15:0] io_SRAM_DQ,
	output        o_SRAM_WE_N,
	output        o_SRAM_CE_N, // no need to handle
	output        o_SRAM_OE_N, // no need to handle
	output        o_SRAM_LB_N, // no need to handle
	output        o_SRAM_UB_N, // no need to handle
	
	// I2C
	input  i_clk_100k,
	output o_I2C_SCLK,
	inout  io_I2C_SDAT,
	
	// AudPlayer
	input  i_AUD_ADCDAT,
	inout  i_AUD_ADCLRCK,
	inout  i_AUD_BCLK,
	inout  i_AUD_DACLRCK,
	output o_AUD_DACDAT

	// SEVENDECODER (optional display)
	// output [5:0] o_record_time,
	// output [5:0] o_play_time,

	// LCD (optional display)
	// input        i_clk_800k,
	// inout  [7:0] o_LCD_DATA,
	// output       o_LCD_EN,
	// output       o_LCD_RS,
	// output       o_LCD_RW,
	// output       o_LCD_ON,
	// output       o_LCD_BLON,

	// LED
	// output  [8:0] o_ledg,
	// output [17:0] o_ledr
);

	// design the FSM and states as you like
	parameter S_I2C        = 0;
	parameter S_IDLE       = 1;
	parameter S_RECD       = 2;
	parameter S_PAUSE      = 3;
	parameter S_PLAY       = 4;

	logic i2c_oen;
	logic [19:0] addr_record, addr_play;
	logic [15:0] data_record, data_play, dac_data;

	assign o_SRAM_ADDR = (state_r == S_RECD) ? addr_record : addr_play[19:0];
	assign io_SRAM_DQ  = (state_r == S_RECD) ? data_record : 16'dz; // sram_dq as output
	assign data_play   = (state_r != S_RECD) ? io_SRAM_DQ : 16'd0; // sram_dq as input
	assign o_SRAM_WE_N = (state_r == S_RECD) ? 1'b0 : 1'b1;

	assign o_SRAM_CE_N = 1'b0;
	assign o_SRAM_OE_N = 1'b0;
	assign o_SRAM_LB_N = 1'b0;
	assign o_SRAM_UB_N = 1'b0;

	// below is a simple example for module division
	// you can design these as you like

	// === I2cInitializer ===
	// sequentially sent out settings to initialize WM8731 with I2C protocal
	I2cInitializer init0(
		.i_rst_n(i_rst_n),
		.i_clk(i_clk_100k),
		.i_start(),
		.o_finished(),
		.o_sclk(o_I2C_SCLK),
		.io_sdat(io_I2C_SDAT),
		.o_oen(i2c_oen) // you are outputing (you are not outputing only when you are "ack"ing.)
	);

	// === AudDSP ===
	// responsible for DSP operations including fast play and slow play at different speed
	// in other words, determine which data addr to be fetch for player 
	AudDSP dsp(
		.i_rst_n(i_rst_n),
		.i_clk(),
		.i_start(),
		.i_pause(),
		.i_speed(), // total 3 bits, use 3 switches
		.i_is_slow(), // 0 for fast play, 1 for slow play, use 1 switch
		.i_slow_mode(), // 0 for constant interpolation, 1 for linear interpolation, use 1 switch
		.i_daclrck(i_AUD_DACLRCK),
		.i_sram_data(data_play),
		.o_dac_data(dac_data),
		.o_sram_addr(addr_play)
	);

	// === AudPlayer ===
	// receive data address from DSP and fetch data to sent to WM8731 with I2S protocal
	AudPlayer player(
		.i_rst_n(i_rst_n),
		.i_bclk(i_AUD_BCLK),
		.i_daclrck(i_AUD_DACLRCK),
		.i_en(), // enable AudPlayer only when playing audio, work with AudDSP
		.i_dac_data(dac_data),
		.o_aud_dacdat(o_AUD_DACDAT)
	);

	// === AudRecorder ===
	// receive data from WM8731 with I2S protocal and save to SRAM
	AudRecorder recorder(
		.i_rst_n(i_rst_n), 
		.i_clk(i_AUD_BCLK),
		.i_lrc(i_AUD_ADCLRCK),
		.i_start(),
		.i_pause(),
		.i_stop(),
		.i_data(i_AUD_ADCDAT),
		.o_address(addr_record),
		.o_data(data_record),
	);

	always @(*) begin
		// design your control here
	end

	always_ff @(posedge i_clk or negedge i_rst_n) begin
		if (!i_rst_n) begin
			
		end
		else begin
			
		end
	end

endmodule
