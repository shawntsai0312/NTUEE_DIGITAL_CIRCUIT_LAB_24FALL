module CoorDecoder(
    input wire i_clk,
    input wire i_rst_n,
    input [10:0] i_H_to_be_rendered,
    input [9:0] i_V_to_be_rendered,
    input signed [10:0] i_x,
    input signed [9:0] i_y,
    output [19:0] o_addr,
);

    

endmodule