module PaddleHandler (
    input i_clk,
    input i_rst_n,
    output o_CS,
    output o_SPC,
    output o_SDI,
    input i_SDO,

    input [7:0] i_level0_lower_bound,
    input [7:0] i_level1_lower_bound,
    input [7:0] i_level2_lower_bound,
    input [7:0] i_level3_lower_bound,
    input [7:0] i_level4_lower_bound,
    input [7:0] i_level5_lower_bound,
    input [7:0] i_level6_lower_bound,
    output [7:0] o_acc_value,
    output reg [2:0] o_level
);
    wire signed [7:0] acc;
    assign o_acc_value = acc;

    ADXL345_ONE_DIR u_ADXL345 (
        .i_clk      (i_clk),
        .i_rst_n    (i_rst_n),
        .o_CS       (o_CS),
        .o_SPC      (o_SPC),
        .o_SDI      (o_SDI),
        .i_SDO      (i_SDO),
        .o_av       (acc)
    );

    always @(*) begin
        o_level = 0;

        if (acc > i_level0_lower_bound) begin
            o_level = 0;
        end else if (acc > i_level1_lower_bound) begin
            o_level = 1;
        end else if (acc > i_level2_lower_bound) begin
            o_level = 2;
        end else if (acc > i_level3_lower_bound) begin
            o_level = 3;
        end else if (acc > i_level4_lower_bound) begin
            o_level = 4;
        end else if (acc > i_level5_lower_bound) begin
            o_level = 5;
        end else if (acc > i_level6_lower_bound) begin
            o_level = 6;
        end else begin
            o_level = 7;
        end
    end

endmodule

module WheelHandler (
    input i_clk,
    input i_rst_n,
    output o_CS,
    output o_SPC,
    output o_SDI,
    input i_SDO,

    input signed [7:0] i_level0_x_bound,
    input signed [7:0] i_level1_x_bound,
    input signed [7:0] i_level2_x_bound,
    input signed [7:0] i_level3_x_bound,
    input signed [7:0] i_level4_x_bound,
    input signed [7:0] i_level5_x_bound,

    output reg signed [3:0] o_level
);
    wire signed [7:0] acc_x, acc_y;
    ADXL345_TWO_DIR u_ADXL345 (
        .i_clk      (i_clk),
        .i_rst_n    (i_rst_n),
        .o_CS       (o_CS),
        .o_SPC      (o_SPC),
        .o_SDI      (o_SDI),
        .i_SDO      (i_SDO),
        .o_av_x     (acc_x),
        .o_av_y     (acc_y)
    );

    always @(*) begin
        o_level = 0;

        if (acc_x >= -i_level0_x_bound && acc_x <= i_level0_x_bound && acc_y <= 0)  o_level = 0;

        if (acc_x >  i_level0_x_bound && acc_x <=  i_level1_x_bound && acc_y <= 0)  o_level = 1;
        if (acc_x >  i_level1_x_bound && acc_x <=  i_level2_x_bound && acc_y <= 0)  o_level = 2;
        if (acc_x >  i_level2_x_bound && acc_x <=  i_level3_x_bound && acc_y <= 0)  o_level = 3;
        if (acc_x >  i_level3_x_bound && acc_x <=  i_level4_x_bound && acc_y <= 0)  o_level = 4;
        if (acc_x >  i_level4_x_bound && acc_x <=  i_level5_x_bound && acc_y <= 0)  o_level = 5;
        if (acc_x >  i_level5_x_bound && acc_y <= 0)  o_level = 6;
        if (acc_x > 0 && acc_y > 0)  o_level = 7;

        if (acc_x < -i_level0_x_bound && acc_x >= -i_level1_x_bound && acc_y <= 0)  o_level = -1;
        if (acc_x < -i_level1_x_bound && acc_x >= -i_level2_x_bound && acc_y <= 0)  o_level = -2;
        if (acc_x < -i_level2_x_bound && acc_x >= -i_level3_x_bound && acc_y <= 0)  o_level = -3;
        if (acc_x < -i_level3_x_bound && acc_x >= -i_level4_x_bound && acc_y <= 0)  o_level = -4;
        if (acc_x < -i_level4_x_bound && acc_x >= -i_level5_x_bound && acc_y <= 0)  o_level = -5;
        if (acc_x < -i_level5_x_bound && acc_y <= 0)  o_level = -6;
        if (acc_x < 0 && acc_y > 0)  o_level = -7;
    end

endmodule