module SramInit(
    input i_clk,
    input i_rst_n,
    input i_start,
    output o_done
);

endmodule