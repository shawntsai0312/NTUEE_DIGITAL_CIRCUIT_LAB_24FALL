module FrameDecoder(
    input i_clk,
    input i_rst_n,


);

endmodule