`timescale 1ns/10ps
`define CYCLE 10.0
`define HCYCLE 5.0
`define MEMFILE "../../tb/AudDSP/golden/mem.txt" // File for SRAM data
`define NUM_MEM_DATA 100
`define SIM_CYCLES 1000000

`define GOLDENFILE "../../tb/AudDSP/golden/linear/linear_7.txt" // File for golden data
`define SPEED 7
`define IS_SLOW 1
`define SLOW_MODE 1
`define NUM_GOLDEN_DATA (`NUM_MEM_DATA * `SPEED)

// `define GOLDENFILE "../../tb/AudDSP/golden/fast/fast_4.txt" // File for golden data
// `define SPEED 4
// `define IS_SLOW 0
// `define SLOW_MODE 1
// `define NUM_GOLDEN_DATA (`NUM_MEM_DATA / `SPEED)    

// `define GOLDENFILE "../../tb/AudDSP/golden/constant/constant_6.txt" // File for golden data
// `define SPEED 6
// `define IS_SLOW 1
// `define SLOW_MODE 0
// `define NUM_GOLDEN_DATA (`NUM_MEM_DATA * `SPEED)

// `define GOLDENFILE "../../tb/AudDSP/golden/normal.txt" // File for golden data
// `define SPEED 1
// `define IS_SLOW 1
// `define SLOW_MODE 0
// `define NUM_GOLDEN_DATA `NUM_MEM_DATA

module tb;
    // Dumping waveform files
    logic i_rst_n, i_clk, i_start, i_pause;
    logic [2:0] i_speed;
    logic i_is_slow, i_slow_mode, i_daclrck;
    logic [15:0] i_sram_data;
    logic [19:0] i_sram_stop_addr;
    logic [15:0] o_dac_data;
    logic o_en;
    logic [19:0] o_sram_addr;

    integer fp_mem, fp_golden;
    // logic [15:0] mem_data [0:`NUM_MEM_DATA-1];
    // logic [15:0] golden_data [0:`NUM_GOLDEN_DATA-1];
    reg [15:0] mem_data[`NUM_MEM_DATA];
    reg [15:0] golden_data[`NUM_GOLDEN_DATA];
    integer i;
    integer error;
    integer diff;

    AudDSP dsp (
        .i_rst_n             (i_rst_n),
        .i_clk               (i_clk),
        .i_start             (i_start),
        // start signal, sent by the controller, not a button press
        .i_pause             (i_pause),
        // pause signal, press to pause, press again to resume
        .i_speed             (i_speed),
        .i_is_slow           (i_is_slow),
        .i_slow_mode         (i_slow_mode),
        .i_daclrck           (i_daclrck),
        // prepare data when low
        .i_sram_data         (i_sram_data),
        .i_sram_stop_addr    (i_sram_stop_addr),
        // the last address to read from SRAM
        .o_dac_data          (o_dac_data),
        .o_en                (o_en),
        // enable signal for AudPlayer, !i_daclrck
        .o_sram_addr         (o_sram_addr)
    );

    // i_clk generation
    initial begin
        i_clk = 1'b1;
    end

    always begin
        #(`HCYCLE) i_clk = ~i_clk;
    end
    
    task load_mem_data;
        input string file_name;
        input integer fp;
        output reg [15:0] data_array[`NUM_MEM_DATA]; // 假設數據是16位寬度
        integer status;
        begin
            fp = $fopen(file_name, "rb");
            if (fp == 0) begin
                $display("Error: Could not open data file.");
                $finish;
            end
            for (integer i = 0; i < `NUM_MEM_DATA; i = i + 1) begin
                status = $fscanf(fp, "%b\n", data_array[i]);
            end
            $fclose(fp);
        end
    endtask

    task load_golden_data;
        input string file_name;
        input integer fp;
        output reg [15:0] data_array[`NUM_GOLDEN_DATA]; // 假設數據是16位寬度
        integer status;
        begin
            fp = $fopen(file_name, "rb");
            if (fp == 0) begin
                $display("Error: Could not open golden data file.");
                $finish;
            end
            for (integer i = 0; i < `NUM_GOLDEN_DATA; i = i + 1) begin
                status = $fscanf(fp, "%b\n", data_array[i]);
            end
            $fclose(fp);
        end
    endtask

    task display_graph_pass;
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;231m░\033[38;5;51;48;5;230m░\033[38;5;109;48;5;247m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;172;48;5;94m░\033[38;5;172;48;5;137m▒\033[38;5;214;48;5;143m▓\033[38;5;80;48;5;254m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;29;48;5;101m▓\033[38;5;208;48;5;173m▒\033[38;5;50;48;5;223m░\033[38;5;138;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[38;5;129;48;5;137m▒\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;166;48;5;180m░\033[38;5;42;48;5;244m▓\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;86;48;5;101m▓\033[38;5;69;48;5;143m▒\033[38;5;179;48;5;136m▒\033[38;5;130;48;5;173m▒\033[38;5;50;48;5;223m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[38;5;80;48;5;101m░\033[38;5;94;48;5;95m▒\033[38;5;130;48;5;52m \033[38;5;180;48;5;94m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;94m░\033[38;5;172;48;5;130m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;43;48;5;223m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;100m▒\033[38;5;172;48;5;94m▒\033[38;5;215;48;5;52m \033[38;5;172;48;5;94m░\033[38;5;179;48;5;173m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;215m░\033[38;5;172;48;5;216m░\033[38;5;179;48;5;186m░\033[38;5;172;48;5;180m▒\033[38;5;50;48;5;224m░\033[38;5;209;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;238m▓\033[38;5;214;48;5;137m▒\033[38;5;172;48;5;94m░\033[38;5;172;48;5;136m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;216m░\033[38;5;214;48;5;186m░\033[38;5;136;48;5;185m░\033[38;5;136;48;5;185m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;223m░\033[38;5;50;48;5;224m░\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;239m▓\033[38;5;69;48;5;180m░\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;172;48;5;58m░\033[38;5;216;48;5;234m \033[38;5;173;48;5;95m▓\033[38;5;208;48;5;137m▓\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;202;48;5;236m▒\033[38;5;208;48;5;95m▓\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;229m \033[38;5;221;48;5;187m▒\033[38;5;87;48;5;230m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;235m▒\033[38;5;50;48;5;187m░\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;95m▒\033[38;5;221;48;5;95m▒\033[38;5;179;48;5;95m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;221m░\033[38;5;94;48;5;221m░\033[38;5;221;48;5;186m░\033[38;5;178;48;5;185m▒\033[38;5;220;48;5;179m▒\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;51;48;5;230m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;203;48;5;186m░\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;222m░\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;137m▓\033[38;5;179;48;5;95m▒\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;144m▓\033[38;5;221;48;5;230m░\033[38;5;94;48;5;224m░\033[38;5;82;48;5;230m░\033[38;5;131;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;50;48;5;180m░\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;101m▓\033[38;5;209;48;5;232m \033[38;5;52;48;5;16m \033[38;5;209;48;5;232m░\033[38;5;208;48;5;237m▓\033[38;5;136;48;5;187m▒\033[38;5;220;48;5;223m▒\033[38;5;29;48;5;224m░\033[38;5;131;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;220;48;5;180m░\033[38;5;178;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;143m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;172;48;5;101m▓\033[38;5;172;48;5;238m▓\033[38;5;208;48;5;235m▓\033[38;5;166;48;5;235m▓\033[38;5;172;48;5;239m▓\033[38;5;136;48;5;144m▓\033[38;5;220;48;5;187m▒\033[38;5;42;48;5;223m▒\033[38;5;174;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;207;48;5;180m░\033[38;5;178;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;95m▒\033[38;5;179;48;5;58m▒\033[38;5;94;48;5;236m░\033[38;5;136;48;5;235m░\033[38;5;220;48;5;235m░\033[38;5;220;48;5;235m░\033[38;5;220;48;5;238m▒\033[38;5;136;48;5;144m▓\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;223m▒\033[38;5;87;48;5;230m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;88;48;5;232m░\033[38;5;50;48;5;187m░\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;223m░\033[38;5;99;48;5;230m▒\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;80;48;5;187m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;51;48;5;230m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;80;48;5;186m░\033[38;5;220;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;94;48;5;223m░\033[38;5;131;48;5;237m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;50;48;5;186m░\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;222m░\033[38;5;214;48;5;223m░\033[38;5;94;48;5;223m░\033[38;5;87;48;5;224m░\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;173;48;5;241m▓\033[38;5;221;48;5;239m▓\033[38;5;43;48;5;180m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;178;48;5;179m▒\033[38;5;220;48;5;179m▒\033[38;5;69;48;5;180m░\033[38;5;50;48;5;187m░\033[38;5;166;48;5;240m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[38;5;130;48;5;242m▓\033[38;5;82;48;5;242m▓\033[38;5;119;48;5;242m▓\033[38;5;65;48;5;242m▓\033[38;5;65;48;5;241m▓\033[38;5;65;48;5;59m▓\033[38;5;191;48;5;59m▓\033[38;5;221;48;5;59m▓\033[38;5;137;48;5;241m▓\033[38;5;202;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[38;5;202;48;5;242m▓\033[38;5;47;48;5;59m▓\033[38;5;50;48;5;187m░\033[38;5;95;48;5;180m▓\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;29;48;5;180m▒\033[38;5;87;48;5;223m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;235m▒\033[38;5;73;48;5;145m▒\033[38;5;51;48;5;230m░\033[38;5;174;48;5;223m▒\033[38;5;221;48;5;223m░\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;84;48;5;180m▒\033[38;5;50;48;5;186m▒\033[38;5;57;48;5;187m▒\033[38;5;51;48;5;187m░\033[38;5;80;48;5;187m░\033[38;5;47;48;5;242m▓\033[38;5;209;48;5;240m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;42;48;5;244m▓\033[38;5;51;48;5;255m░\033[38;5;50;48;5;224m▒\033[38;5;94;48;5;187m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;173m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;179;48;5;180m▒\033[38;5;50;48;5;187m░\033[38;5;29;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;87;48;5;255m░\033[38;5;29;48;5;224m░\033[38;5;172;48;5;223m░\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;143m▒\033[38;5;68;48;5;180m▒\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;248m▒\033[38;5;214;48;5;224m░\033[38;5;214;48;5;186m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;51;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;51;48;5;255m░\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;143m▒\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;220;48;5;143m▒\033[38;5;51;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;255m░\033[38;5;172;48;5;187m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;178;48;5;143m▒\033[38;5;80;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;236m▒\033[38;5;69;48;5;223m░\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;172;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;178;48;5;179m▒\033[38;5;42;48;5;179m▒\033[38;5;36;48;5;101m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;236m▒\033[38;5;185;48;5;187m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;163;48;5;180m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;235m▒\033[38;5;130;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;32;48;5;179m▒\033[38;5;47;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;224m░\033[38;5;179;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;67;48;5;179m▒\033[38;5;78;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;50;48;5;223m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;25;48;5;179m▒\033[38;5;72;48;5;101m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m▒\033[38;5;179;48;5;223m░\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;67;48;5;180m▒\033[38;5;130;48;5;241m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;93;48;5;223m░\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;173m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;118;48;5;223m▒\033[38;5;84;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;45;48;5;223m░\033[38;5;136;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;237m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;233m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;235m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;240m▒\033[38;5;94;48;5;101m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;234m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;45;48;5;186m▒\033[38;5;65;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;99;48;5;187m▓\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;242;48;5;241m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;232;48;5;232m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;252;48;5;252m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;232m \033[38;5;221;48;5;101m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;234;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;57;48;5;180m░\033[38;5;113;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;51;48;5;187m░\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;236m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;234;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;250;48;5;250m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;248;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;236m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;50;48;5;186m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;245;48;5;245m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;236;48;5;236m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;249;48;5;249m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;241;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;237;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;249;48;5;249m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;50;48;5;223m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;223m░\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;75;48;5;180m░\033[38;5;50;48;5;222m░\033[38;5;35;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;245;48;5;245m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;247;48;5;247m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;235;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;235;48;5;235m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;239;48;5;239m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;242;48;5;241m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;130;48;5;232m \033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;31;48;5;179m░\033[38;5;78;48;5;101m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[38;5;86;48;5;138m▓\033[38;5;50;48;5;186m░\033[38;5;136;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;209;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;237;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;246;48;5;246m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;235m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;232;48;5;232m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;234;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;230;48;5;180m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;47;48;5;180m▒\033[38;5;202;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;249m▒\033[38;5;62;48;5;186m░\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;209;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;245;48;5;245m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;234;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;240;48;5;240m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;249;48;5;249m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;251;48;5;251m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;234;48;5;234m▓\033[38;5;233;48;5;233m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;237;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;172;48;5;95m▓\033[38;5;49;48;5;187m▒\033[38;5;208;48;5;223m░\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;179m▒\033[38;5;130;48;5;173m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;42;48;5;95m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;204;48;5;180m▓\033[38;5;220;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;32;48;5;186m▒\033[38;5;87;48;5;229m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;144m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;216;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;242;48;5;242m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;232;48;5;232m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;252;48;5;252m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;234;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;50;48;5;187m░\033[38;5;1;48;5;232m░\033[0m \033[38;5;50;48;5;252m▒\033[38;5;190;48;5;187m░\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;165;48;5;180m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;223m░\033[38;5;136;48;5;144m▒\033[38;5;178;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;179m▒\033[38;5;50;48;5;187m░\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[38;5;51;48;5;223m░\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;233m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;202;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;209;48;5;16m \033[38;5;94;48;5;179m▒\033[38;5;214;48;5;95m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;239m▓\033[38;5;35;48;5;187m░\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[38;5;123;48;5;230m░\033[38;5;26;48;5;186m░\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;200;48;5;180m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;50;48;5;180m░\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;50;48;5;187m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;224m░\033[38;5;214;48;5;144m▓\033[38;5;214;48;5;137m▓\033[38;5;94;48;5;233m▒\033[38;5;202;48;5;16m \033[38;5;202;48;5;16m \033[38;5;166;48;5;16m \033[38;5;94;48;5;232m░\033[38;5;94;48;5;137m▓\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;143m▒\033[38;5;94;48;5;233m▒\033[38;5;166;48;5;232m \033[38;5;202;48;5;16m \033[38;5;209;48;5;16m \033[38;5;214;48;5;234m░\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;58m▒\033[38;5;202;48;5;16m \033[38;5;209;48;5;16m \033[38;5;209;48;5;16m \033[38;5;166;48;5;232m \033[38;5;94;48;5;239m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;236m▒\033[38;5;172;48;5;232m \033[38;5;216;48;5;16m \033[38;5;222;48;5;232m \033[38;5;221;48;5;235m▒\033[38;5;221;48;5;95m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;237m▒\033[38;5;222;48;5;233m░\033[38;5;209;48;5;16m \033[38;5;172;48;5;232m \033[38;5;179;48;5;236m▒\033[38;5;214;48;5;101m▓\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;77;48;5;180m▒\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;191;48;5;180m░\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;156;48;5;180m░\033[38;5;84;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;88;48;5;232m░\033[38;5;71;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;51;48;5;223m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;181m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;179;48;5;180m░\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;50;48;5;223m░\033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;45;48;5;180m░\033[38;5;84;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;88;48;5;232m░\033[38;5;69;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;47;48;5;186m░\033[38;5;166;48;5;240m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;144m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;179;48;5;180m░\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;167;48;5;232m░\033[0m \033[0m \033[0m \033[38;5;87;48;5;223m░\033[38;5;220;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;80;48;5;180m░\033[38;5;84;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;88;48;5;232m░\033[38;5;29;48;5;180m▓\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;214;48;5;186m▒\033[38;5;50;48;5;224m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;93;48;5;186m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m░\033[38;5;178;48;5;186m░\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;87;48;5;230m░\033[0m \033[0m \033[0m \033[38;5;47;48;5;186m▒\033[38;5;221;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;45;48;5;180m░\033[38;5;84;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;50;48;5;181m░\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;186m▒\033[38;5;50;48;5;224m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;50;48;5;223m░\033[0m \033[0m \033[38;5;50;48;5;253m░\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;45;48;5;180m▒\033[38;5;84;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;144m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;99;48;5;186m▒\033[38;5;131;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;223m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;50;48;5;223m░\033[0m \033[0m \033[38;5;80;48;5;187m░\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;31;48;5;180m▓\033[38;5;209;48;5;240m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;178;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;87;48;5;229m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;51;48;5;187m░\033[38;5;88;48;5;232m░\033[0m \033[38;5;80;48;5;253m░\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;50;48;5;180m░\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;223m░\033[38;5;87;48;5;230m░\033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;221;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;144m▒\033[38;5;86;48;5;101m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;88;48;5;232m░\033[38;5;50;48;5;186m░\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;50;48;5;224m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;50;48;5;223m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;99;48;5;180m░\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;206;48;5;180m░\033[38;5;138;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m░\033[38;5;178;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;137m▓\033[38;5;80;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;223m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;185m░\033[38;5;50;48;5;223m░\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;102m▓\033[38;5;178;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;29;48;5;101m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;109;48;5;245m▓\033[38;5;220;48;5;143m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;137m▒\033[38;5;80;48;5;186m░\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;252m▒\033[38;5;78;48;5;187m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;50;48;5;223m░\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;95;48;5;240m▓\033[38;5;44;48;5;180m░\033[38;5;221;48;5;137m▓\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;220;48;5;180m▒\033[38;5;116;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;50;48;5;144m░\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;220;48;5;137m▒\033[38;5;220;48;5;137m▒\033[38;5;220;48;5;137m▒\033[38;5;80;48;5;187m░\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;251m▒\033[38;5;214;48;5;180m▒\033[38;5;220;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;52;48;5;180m░\033[38;5;103;48;5;186m▓\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;186m░\033[38;5;178;48;5;143m▓\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;43;48;5;180m░\033[38;5;43;48;5;102m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;101m▓\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;62;48;5;101m░\033[38;5;29;48;5;243m▓\033[0m \033[0m \033[0m \033[38;5;202;48;5;241m▓\033[38;5;86;48;5;179m▒\033[38;5;220;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;50;48;5;186m░\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[38;5;174;48;5;236m▒\033[38;5;50;48;5;186m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;50;48;5;180m░\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[38;5;209;48;5;239m▓\033[38;5;44;48;5;144m░\033[38;5;178;48;5;143m▓\033[38;5;136;48;5;143m▓\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;187m▒\033[38;5;44;48;5;187m░\033[38;5;138;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▓\033[38;5;161;48;5;187m░\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;220;48;5;143m▒\033[38;5;136;48;5;143m▓\033[38;5;179;48;5;137m▒\033[38;5;130;48;5;137m▓\033[38;5;42;48;5;243m▓\033[0m \033[0m \033[0m \033[38;5;50;48;5;187m▒\033[38;5;220;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;78;48;5;242m▓\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;69;48;5;179m░\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[38;5;116;48;5;144m▒\033[38;5;136;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;187m▒\033[38;5;50;48;5;250m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;51;48;5;230m░\033[38;5;94;48;5;187m▒\033[38;5;214;48;5;187m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;214;48;5;137m▒\033[38;5;39;48;5;101m▒\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[38;5;80;48;5;187m▒\033[38;5;178;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;114;48;5;179m▒\033[38;5;116;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[38;5;116;48;5;249m▒\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;209;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;224m░\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;86;48;5;137m▒\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;178;48;5;179m▒\033[38;5;80;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m░\033[38;5;214;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;50;48;5;180m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[38;5;50;48;5;245m▒\033[38;5;214;48;5;101m▓\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;84;48;5;187m▒\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;239m▓\033[38;5;33;48;5;187m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;101m▒\033[38;5;221;48;5;58m▒\033[38;5;94;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;50;48;5;138m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;82;48;5;180m░\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;42;48;5;241m▓\033[38;5;179;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;27;48;5;179m░\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[38;5;138;48;5;239m▓\033[38;5;85;48;5;137m░\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m░\033[38;5;214;48;5;186m░\033[38;5;214;48;5;186m░\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;47;48;5;187m░\033[38;5;50;48;5;249m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;51;48;5;187m░\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m░\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m░\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;144m▓\033[38;5;50;48;5;180m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;180m░\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;47;48;5;243m▓\033[38;5;57;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;173m▒\033[38;5;36;48;5;223m░\033[0m \033[0m \033[0m \033[0m \033[38;5;116;48;5;249m▒\033[38;5;136;48;5;95m▓\033[38;5;221;48;5;95m▒\033[38;5;94;48;5;94m▒\033[38;5;214;48;5;101m▒\033[38;5;214;48;5;144m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m░\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;199;48;5;187m▒\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;51;48;5;223m░\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;187m▒\033[38;5;221;48;5;223m░\033[38;5;221;48;5;187m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;221;48;5;144m▓\033[38;5;80;48;5;254m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;238m▓\033[38;5;40;48;5;179m░\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;80;48;5;186m░\033[38;5;131;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;238m▓\033[38;5;200;48;5;186m▓\033[38;5;214;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;208;48;5;180m▓\033[38;5;174;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▓\033[38;5;32;48;5;137m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;178;48;5;222m░\033[38;5;220;48;5;180m▒\033[38;5;220;48;5;180m▒\033[38;5;80;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;246m▓\033[38;5;77;48;5;138m░\033[38;5;136;48;5;144m▓\033[38;5;83;48;5;223m░\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;220;48;5;180m▒\033[38;5;69;48;5;180m░\033[38;5;80;48;5;253m░\033[38;5;209;48;5;236m▓\033[38;5;80;48;5;253m░\033[38;5;131;48;5;237m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;84;48;5;180m░\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;136;48;5;143m▒\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;50;48;5;180m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m░\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;50;48;5;223m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m▒\033[38;5;220;48;5;144m▓\033[38;5;178;48;5;144m▓\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;187m▒\033[38;5;94;48;5;186m▒\033[38;5;136;48;5;187m▒\033[38;5;27;48;5;187m░\033[38;5;119;48;5;101m░\033[38;5;116;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;131;48;5;237m▓\033[38;5;131;48;5;237m▓\033[38;5;87;48;5;255m░\033[38;5;87;48;5;254m░\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;149;48;5;243m▓\033[38;5;101;48;5;187m▓\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;162;48;5;180m▒\033[38;5;174;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[0m \033[38;5;131;48;5;237m▓\033[38;5;80;48;5;187m░\033[38;5;86;48;5;187m░\033[38;5;220;48;5;187m░\033[38;5;80;48;5;253m░\033[38;5;131;48;5;237m▓\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;185;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;101;48;5;243m▓\033[38;5;156;48;5;180m░\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;50;48;5;180m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;123;48;5;230m░\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;62;48;5;180m░\033[38;5;167;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;137;48;5;243m▓\033[38;5;192;48;5;181m░\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;50;48;5;181m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;211;48;5;187m░\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;220;48;5;179m▒\033[38;5;220;48;5;143m▒\033[38;5;50;48;5;187m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;204;48;5;180m░\033[38;5;221;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;69;48;5;143m░\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m░\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;144m▒\033[38;5;87;48;5;224m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;161;48;5;143m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;244m▓\033[38;5;35;48;5;180m░\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;50;48;5;180m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;224m░\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;40;48;5;180m░\033[38;5;50;48;5;253m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;45;48;5;241m▓\033[38;5;25;48;5;138m░\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;144m▒\033[38;5;221;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;143;48;5;180m▒\033[38;5;93;48;5;150m▒\033[38;5;80;48;5;187m░\033[38;5;116;48;5;250m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;224m░\033[38;5;178;48;5;144m▓\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;51;48;5;143m░\033[38;5;45;48;5;143m░\033[38;5;80;48;5;143m▒\033[38;5;45;48;5;144m░\033[38;5;50;48;5;145m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;88;48;5;232m░\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m");
    endtask

    task display_graph_fail;
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;88;48;5;232m░\033[38;5;116;48;5;250m▒\033[38;5;62;48;5;101m▒\033[38;5;220;48;5;240m▓\033[38;5;178;48;5;95m▓\033[38;5;69;48;5;101m░\033[38;5;44;48;5;144m░\033[38;5;80;48;5;253m░\033[38;5;87;48;5;230m░\033[38;5;87;48;5;230m░\033[38;5;87;48;5;230m░\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;239m▓\033[38;5;52;48;5;101m░\033[38;5;221;48;5;94m▒\033[38;5;94;48;5;94m▒\033[38;5;214;48;5;94m▒\033[38;5;179;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;101m▓\033[38;5;172;48;5;101m▓\033[38;5;172;48;5;101m▓\033[38;5;130;48;5;101m▓\033[38;5;172;48;5;137m▓\033[38;5;130;48;5;137m▓\033[38;5;172;48;5;137m▓\033[38;5;32;48;5;137m░\033[38;5;26;48;5;137m░\033[38;5;148;48;5;137m▒\033[38;5;209;48;5;144m░\033[38;5;50;48;5;144m░\033[38;5;50;48;5;187m░\033[38;5;50;48;5;187m░\033[38;5;116;48;5;181m▒\033[38;5;35;48;5;242m▓\033[38;5;47;48;5;243m▓\033[38;5;166;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;39;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;94m▒\033[38;5;208;48;5;240m▒\033[38;5;36;48;5;101m░\033[38;5;86;48;5;246m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;224m░\033[38;5;50;48;5;180m░\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;130;48;5;58m \033[38;5;130;48;5;58m░\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;95m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;58m▒\033[38;5;130;48;5;236m▒\033[38;5;50;48;5;101m░\033[38;5;50;48;5;245m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;238m▓\033[38;5;50;48;5;187m░\033[38;5;179;48;5;143m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;58m░\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;58m \033[38;5;172;48;5;235m \033[38;5;172;48;5;58m▒\033[38;5;50;48;5;101m░\033[38;5;47;48;5;241m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;236m▒\033[38;5;80;48;5;181m░\033[38;5;179;48;5;144m▓\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;95m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;52m \033[38;5;215;48;5;52m \033[38;5;208;48;5;58m░\033[38;5;180;48;5;239m▒\033[38;5;43;48;5;138m▒\033[38;5;49;48;5;245m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m▒\033[38;5;220;48;5;137m▓\033[38;5;172;48;5;144m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;94m░\033[38;5;172;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;130m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;137;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;215;48;5;52m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m▒\033[38;5;57;48;5;95m▓\033[38;5;50;48;5;181m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;245m▓\033[38;5;50;48;5;101m▓\033[38;5;220;48;5;59m▓\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;173m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;95m▒\033[38;5;215;48;5;58m░\033[38;5;202;48;5;52m \033[38;5;216;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m▒\033[38;5;166;48;5;58m▒\033[38;5;69;48;5;95m▒\033[38;5;50;48;5;181m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;116;48;5;248m▒\033[38;5;190;48;5;234m▒\033[38;5;58;48;5;234m \033[38;5;172;48;5;95m▒\033[38;5;130;48;5;173m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;130m░\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;95m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;130m▒\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;52m \033[38;5;216;48;5;52m \033[38;5;216;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;95m▒\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;246m▒\033[38;5;190;48;5;237m▓\033[38;5;136;48;5;238m▓\033[38;5;137;48;5;95m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;130m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;58m▒\033[38;5;76;48;5;238m▓\033[38;5;74;48;5;237m▓\033[38;5;110;48;5;233m▒\033[38;5;137;48;5;232m▓\033[38;5;202;48;5;232m \033[38;5;209;48;5;232m \033[38;5;52;48;5;233m \033[38;5;202;48;5;52m \033[38;5;208;48;5;94m▒\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;137m▒\033[38;5;180;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;130m░\033[38;5;166;48;5;130m░\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;1m░\033[38;5;202;48;5;52m \033[38;5;202;48;5;52m \033[38;5;216;48;5;52m \033[38;5;202;48;5;52m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;172;48;5;58m▒\033[38;5;21;48;5;95m░\033[38;5;73;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;101m░\033[38;5;179;48;5;240m▒\033[38;5;179;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;173;48;5;58m▒\033[38;5;209;48;5;52m▒\033[38;5;204;48;5;239m▓\033[38;5;60;48;5;60m▓\033[38;5;68;48;5;67m▓\033[38;5;26;48;5;66m▓\033[38;5;26;48;5;241m▓\033[38;5;209;48;5;59m▓\033[38;5;166;48;5;95m▓\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;172;48;5;180m░\033[38;5;130;48;5;180m░\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;130m░\033[38;5;180;48;5;130m░\033[38;5;180;48;5;130m░\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;27;48;5;101m▒\033[38;5;80;48;5;253m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;50;48;5;181m▒\033[38;5;121;48;5;240m░\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;208;48;5;94m░\033[38;5;172;48;5;101m▒\033[38;5;220;48;5;101m▓\033[38;5;74;48;5;245m▓\033[38;5;208;48;5;248m▓\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;179;48;5;239m▒\033[38;5;176;48;5;101m▒\033[38;5;137;48;5;59m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;50;48;5;250m▒\033[38;5;94;48;5;101m░\033[38;5;172;48;5;238m▓\033[38;5;172;48;5;236m▒\033[38;5;172;48;5;235m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;131m▒\033[38;5;172;48;5;137m▒\033[38;5;220;48;5;144m▓\033[38;5;25;48;5;246m▓\033[38;5;45;48;5;246m▓\033[38;5;144;48;5;144m▓\033[38;5;220;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;187m▒\033[38;5;214;48;5;187m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;130m▒\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;172;48;5;58m▒\033[38;5;179;48;5;238m▒\033[38;5;21;48;5;59m░\033[38;5;50;48;5;138m▒\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;238m▓\033[38;5;80;48;5;102m░\033[38;5;220;48;5;238m▓\033[38;5;220;48;5;235m▒\033[38;5;220;48;5;235m▒\033[38;5;178;48;5;234m░\033[38;5;214;48;5;235m░\033[38;5;179;48;5;58m░\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;94;48;5;144m▓\033[38;5;39;48;5;109m▓\033[38;5;25;48;5;67m▓\033[38;5;35;48;5;248m▓\033[38;5;112;48;5;151m▓\033[38;5;190;48;5;187m▓\033[38;5;144;48;5;187m▓\033[38;5;178;48;5;187m▓\033[38;5;178;48;5;187m▓\033[38;5;214;48;5;188m▓\033[38;5;179;48;5;188m▒\033[38;5;172;48;5;187m▒\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;95m▓\033[38;5;50;48;5;181m░\033[38;5;86;48;5;246m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;145m▓\033[38;5;216;48;5;239m░\033[38;5;58;48;5;232m \033[38;5;58;48;5;232m \033[38;5;58;48;5;233m \033[38;5;58;48;5;233m \033[38;5;220;48;5;233m \033[38;5;136;48;5;235m░\033[38;5;221;48;5;58m▒\033[38;5;179;48;5;95m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;101m▒\033[38;5;214;48;5;101m▒\033[38;5;94;48;5;137m▒\033[38;5;112;48;5;244m▓\033[38;5;39;48;5;60m▓\033[38;5;35;48;5;245m▓\033[38;5;190;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;172;48;5;181m▓\033[38;5;179;48;5;187m▓\033[38;5;130;48;5;187m▒\033[38;5;130;48;5;187m▒\033[38;5;130;48;5;187m▒\033[38;5;172;48;5;187m▒\033[38;5;172;48;5;187m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;95m▓\033[38;5;80;48;5;181m▒\033[38;5;43;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;131;48;5;240m▓\033[38;5;143;48;5;232m▒\033[38;5;58;48;5;232m \033[38;5;190;48;5;232m \033[38;5;220;48;5;232m \033[38;5;136;48;5;232m \033[38;5;222;48;5;232m \033[38;5;172;48;5;233m \033[38;5;221;48;5;235m░\033[38;5;94;48;5;240m▒\033[38;5;214;48;5;101m▓\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;214;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;221;48;5;94m▒\033[38;5;220;48;5;58m▒\033[38;5;143;48;5;237m▒\033[38;5;178;48;5;239m▓\033[38;5;221;48;5;95m▓\033[38;5;179;48;5;137m▓\033[38;5;214;48;5;144m▓\033[38;5;136;48;5;144m▓\033[38;5;221;48;5;144m▒\033[38;5;221;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;221;48;5;58m▒\033[38;5;221;48;5;95m▓\033[38;5;50;48;5;144m░\033[38;5;149;48;5;59m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;116;48;5;246m▒\033[38;5;190;48;5;233m▓\033[38;5;155;48;5;16m \033[38;5;58;48;5;232m \033[38;5;220;48;5;232m \033[38;5;136;48;5;232m \033[38;5;214;48;5;232m \033[38;5;136;48;5;234m░\033[38;5;221;48;5;238m▒\033[38;5;94;48;5;95m▓\033[38;5;179;48;5;101m▓\033[38;5;214;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;94m▒\033[38;5;221;48;5;58m▒\033[38;5;178;48;5;58m░\033[38;5;172;48;5;234m \033[38;5;172;48;5;233m \033[38;5;221;48;5;58m░\033[38;5;221;48;5;95m▒\033[38;5;221;48;5;101m▓\033[38;5;94;48;5;143m▓\033[38;5;221;48;5;144m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;143m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;131m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;179;48;5;94m▒\033[38;5;214;48;5;94m▒\033[38;5;94;48;5;94m▒\033[38;5;94;48;5;95m▒\033[38;5;50;48;5;144m░\033[38;5;49;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;241;48;5;240m▓\033[38;5;80;48;5;242m▒\033[38;5;143;48;5;235m▓\033[38;5;220;48;5;235m▒\033[38;5;220;48;5;235m▒\033[38;5;220;48;5;235m▒\033[38;5;178;48;5;236m▒\033[38;5;221;48;5;238m▓\033[38;5;94;48;5;59m▓\033[38;5;214;48;5;95m▓\033[38;5;214;48;5;95m▒\033[38;5;94;48;5;58m▒\033[38;5;221;48;5;58m▒\033[38;5;221;48;5;58m▒\033[38;5;221;48;5;58m░\033[38;5;222;48;5;234m \033[38;5;94;48;5;234m \033[38;5;136;48;5;58m░\033[38;5;221;48;5;58m▒\033[38;5;136;48;5;95m▒\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;137m▓\033[38;5;94;48;5;144m▓\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;131m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;214;48;5;94m▒\033[38;5;221;48;5;94m▒\033[38;5;221;48;5;95m▒\033[38;5;80;48;5;181m▒\033[38;5;50;48;5;246m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;109;48;5;248m▓\033[38;5;66;48;5;244m▓\033[38;5;109;48;5;241m▓\033[38;5;116;48;5;243m▒\033[38;5;80;48;5;243m▒\033[38;5;220;48;5;59m▒\033[38;5;136;48;5;238m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;58m░\033[38;5;136;48;5;58m▒\033[38;5;136;48;5;240m▒\033[38;5;136;48;5;101m▒\033[38;5;221;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;137m▓\033[38;5;136;48;5;143m▓\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;131m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;179;48;5;94m▒\033[38;5;94;48;5;94m▒\033[38;5;136;48;5;94m▒\033[38;5;178;48;5;94m▒\033[38;5;33;48;5;101m▒\033[38;5;80;48;5;187m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[38;5;80;48;5;144m▒\033[38;5;220;48;5;101m▓\033[38;5;178;48;5;101m▓\033[38;5;178;48;5;101m▒\033[38;5;136;48;5;95m▒\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;101m▓\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;143m▓\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;216;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;179;48;5;94m▒\033[38;5;214;48;5;95m▒\033[38;5;50;48;5;144m░\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m▒\033[38;5;220;48;5;101m▓\033[38;5;178;48;5;101m▓\033[38;5;221;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;214;48;5;137m▓\033[38;5;214;48;5;137m▓\033[38;5;179;48;5;144m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;216;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;215;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;130;48;5;95m▒\033[38;5;55;48;5;138m▒\033[38;5;50;48;5;144m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;252m▒\033[38;5;220;48;5;144m▓\033[38;5;136;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;131m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;166;48;5;94m▒\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m▒\033[38;5;130;48;5;95m▒\033[38;5;84;48;5;138m▒\033[38;5;86;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;252m▒\033[38;5;178;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;130;48;5;144m▓\033[38;5;130;48;5;144m▓\033[38;5;130;48;5;144m▓\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;144m▒\033[38;5;179;48;5;144m▒\033[38;5;221;48;5;144m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;95m▒\033[38;5;226;48;5;144m░\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;252m▒\033[38;5;214;48;5;249m▓\033[38;5;172;48;5;180m▓\033[38;5;172;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▓\033[38;5;130;48;5;180m▓\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;144m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;180;48;5;130m░\033[38;5;180;48;5;130m░\033[38;5;166;48;5;130m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;173;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;208;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;202;48;5;52m░\033[38;5;166;48;5;58m░\033[38;5;180;48;5;94m░\033[38;5;208;48;5;94m▒\033[38;5;172;48;5;95m▓\033[38;5;80;48;5;144m░\033[38;5;131;48;5;237m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;252m▒\033[38;5;172;48;5;249m▓\033[38;5;172;48;5;95m▓\033[38;5;130;48;5;234m▓\033[38;5;130;48;5;234m▓\033[38;5;130;48;5;234m▓\033[38;5;172;48;5;234m▓\033[38;5;130;48;5;234m▓\033[38;5;130;48;5;234m▓\033[38;5;172;48;5;234m▓\033[38;5;172;48;5;234m▓\033[38;5;130;48;5;234m▓\033[38;5;130;48;5;234m▓\033[38;5;214;48;5;234m▓\033[38;5;94;48;5;234m▒\033[38;5;221;48;5;233m▒\033[38;5;222;48;5;233m░\033[38;5;179;48;5;236m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;58m░\033[38;5;209;48;5;232m \033[38;5;209;48;5;232m \033[38;5;209;48;5;232m \033[38;5;209;48;5;232m \033[38;5;209;48;5;232m \033[38;5;202;48;5;233m \033[38;5;180;48;5;94m░\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;234m░\033[38;5;216;48;5;232m \033[38;5;216;48;5;232m \033[38;5;202;48;5;233m \033[38;5;202;48;5;232m \033[38;5;215;48;5;234m░\033[38;5;180;48;5;58m▒\033[38;5;208;48;5;234m░\033[38;5;202;48;5;232m \033[38;5;216;48;5;232m \033[38;5;209;48;5;232m \033[38;5;216;48;5;232m \033[38;5;130;48;5;234m░\033[38;5;208;48;5;58m░\033[38;5;208;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;202;48;5;52m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;130;48;5;95m▒\033[38;5;43;48;5;101m░\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;116;48;5;246m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;137m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;215;48;5;52m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;50;48;5;180m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;238;48;5;238m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;172;48;5;236m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;234m \033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;52m░\033[38;5;166;48;5;52m░\033[38;5;166;48;5;52m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;62;48;5;101m▒\033[38;5;50;48;5;144m▓\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;238m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;235;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;253;48;5;253m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;234m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;52m░\033[38;5;202;48;5;52m \033[38;5;202;48;5;52m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;58m▒\033[38;5;201;48;5;101m░\033[38;5;29;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;238m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;252m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;249;48;5;249m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;234m░\033[38;5;166;48;5;94m▒\033[38;5;202;48;5;58m░\033[38;5;202;48;5;52m░\033[38;5;216;48;5;52m \033[38;5;216;48;5;52m \033[38;5;166;48;5;52m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m▒\033[38;5;50;48;5;144m▒\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;238m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;248;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;237;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;235m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;52m░\033[38;5;216;48;5;52m \033[38;5;216;48;5;52m \033[38;5;166;48;5;52m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;52m░\033[38;5;179;48;5;236m▒\033[38;5;80;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;237m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;234;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;235;48;5;235m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;232;48;5;232m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;238;48;5;238m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;234m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;52m░\033[38;5;202;48;5;52m \033[38;5;202;48;5;52m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;208;48;5;52m \033[38;5;130;48;5;234m░\033[38;5;190;48;5;239m░\033[38;5;109;48;5;248m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;243;48;5;243m▓\033[38;5;73;48;5;237m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;7;48;5;7m▓\033[38;5;7;48;5;7m▓\033[38;5;251;48;5;251m▓\033[38;5;7;48;5;7m▓\033[38;5;7;48;5;7m▓\033[38;5;7;48;5;7m▓\033[38;5;251;48;5;251m▓\033[38;5;7;48;5;7m▓\033[38;5;232;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;252;48;5;252m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;209;48;5;232m \033[38;5;202;48;5;52m \033[38;5;216;48;5;234m \033[38;5;216;48;5;234m \033[38;5;202;48;5;52m \033[38;5;166;48;5;52m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;215;48;5;52m \033[38;5;208;48;5;235m░\033[38;5;130;48;5;234m░\033[38;5;50;48;5;243m▒\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;237m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;249;48;5;249m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;16m \033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;215;48;5;58m░\033[38;5;215;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;215;48;5;52m░\033[38;5;84;48;5;236m▒\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;243;48;5;242m▓\033[38;5;50;48;5;237m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;237m▓\033[38;5;179;48;5;240m▓\033[38;5;172;48;5;236m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;242;48;5;241m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;233;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;239;48;5;239m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;233;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;243;48;5;242m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;52m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;215;48;5;52m \033[38;5;208;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;172;48;5;101m▓\033[38;5;179;48;5;144m▓\033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;235m▒\033[38;5;94;48;5;233m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;248;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;252;48;5;252m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;7;48;5;7m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;234m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;52m░\033[38;5;166;48;5;52m \033[38;5;215;48;5;52m░\033[38;5;215;48;5;52m░\033[38;5;215;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;240m▒\033[38;5;50;48;5;101m░\033[38;5;47;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;245m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;232m \033[38;5;179;48;5;144m▓\033[38;5;179;48;5;144m▒\033[38;5;179;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;238m▓\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;233m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;45;48;5;240m▒\033[38;5;202;48;5;241m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;253m░\033[38;5;76;48;5;144m░\033[38;5;221;48;5;237m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;232m \033[38;5;136;48;5;101m▓\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;144m▓\033[38;5;179;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;237m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;16m \033[38;5;215;48;5;233m \033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;16m \033[38;5;215;48;5;52m░\033[38;5;180;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;45;48;5;238m░\033[38;5;209;48;5;59m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;162;48;5;144m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m▒\033[38;5;38;48;5;240m▒\033[38;5;202;48;5;241m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;70;48;5;143m░\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;50;48;5;101m▒\033[38;5;174;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;55;48;5;137m▓\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;143m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;208;48;5;237m▒\033[38;5;69;48;5;239m░\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;76;48;5;137m░\033[38;5;221;48;5;101m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m \033[38;5;130;48;5;58m░\033[38;5;130;48;5;52m░\033[38;5;130;48;5;236m░\033[38;5;130;48;5;236m▒\033[38;5;209;48;5;240m▒\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;119;48;5;137m░\033[38;5;221;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;215;48;5;52m \033[38;5;215;48;5;52m \033[38;5;130;48;5;52m \033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;130;48;5;237m▒\033[38;5;82;48;5;238m▒\033[38;5;49;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;46;48;5;137m░\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;215;48;5;52m \033[38;5;215;48;5;52m \033[38;5;215;48;5;52m \033[38;5;130;48;5;52m \033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;58m▒\033[38;5;77;48;5;238m▒\033[38;5;50;48;5;247m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;46;48;5;137m░\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;95m▒\033[38;5;214;48;5;94m▒\033[38;5;94;48;5;94m▒\033[38;5;94;48;5;94m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;52m \033[38;5;215;48;5;52m \033[38;5;166;48;5;234m \033[38;5;215;48;5;52m \033[38;5;208;48;5;52m \033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;58m▒\033[38;5;70;48;5;95m░\033[38;5;50;48;5;181m▒\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;253m░\033[38;5;32;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;94m▒\033[38;5;214;48;5;58m░\033[38;5;214;48;5;58m \033[38;5;214;48;5;58m \033[38;5;94;48;5;58m▒\033[38;5;94;48;5;95m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;94m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;130m▒\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;215;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;52m \033[38;5;215;48;5;234m \033[38;5;166;48;5;234m \033[38;5;166;48;5;234m \033[38;5;215;48;5;52m \033[38;5;130;48;5;52m \033[38;5;130;48;5;52m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;104;48;5;95m▒\033[38;5;42;48;5;101m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;239m▓\033[38;5;109;48;5;247m▓\033[38;5;80;48;5;187m░\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;95m▒\033[38;5;136;48;5;58m▒\033[38;5;221;48;5;58m \033[38;5;214;48;5;235m \033[38;5;222;48;5;235m \033[38;5;214;48;5;58m \033[38;5;94;48;5;58m░\033[38;5;214;48;5;94m▒\033[38;5;214;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;130;48;5;58m░\033[38;5;172;48;5;52m \033[38;5;215;48;5;234m \033[38;5;166;48;5;233m \033[38;5;166;48;5;234m \033[38;5;215;48;5;234m \033[38;5;130;48;5;52m \033[38;5;172;48;5;52m░\033[38;5;172;48;5;58m░\033[38;5;222;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;236m▒\033[38;5;36;48;5;95m▒\033[38;5;174;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;109;48;5;247m▓\033[38;5;109;48;5;246m▓\033[38;5;80;48;5;188m░\033[38;5;208;48;5;250m▒\033[38;5;101;48;5;144m▓\033[38;5;144;48;5;143m▓\033[38;5;220;48;5;143m▓\033[38;5;221;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;178;48;5;101m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;58m░\033[38;5;178;48;5;58m░\033[38;5;221;48;5;58m░\033[38;5;94;48;5;58m░\033[38;5;214;48;5;58m░\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;173m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;52m \033[38;5;166;48;5;234m \033[38;5;166;48;5;233m \033[38;5;130;48;5;234m \033[38;5;172;48;5;234m \033[38;5;222;48;5;235m \033[38;5;222;48;5;235m \033[38;5;214;48;5;235m \033[38;5;214;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;222;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;56;48;5;238m░\033[38;5;72;48;5;59m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;80;48;5;187m░\033[38;5;44;48;5;187m░\033[38;5;29;48;5;144m░\033[38;5;144;48;5;101m▓\033[38;5;144;48;5;101m▓\033[38;5;144;48;5;101m▓\033[38;5;143;48;5;101m▓\033[38;5;143;48;5;101m▓\033[38;5;143;48;5;101m▓\033[38;5;220;48;5;101m▒\033[38;5;220;48;5;101m▒\033[38;5;136;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;137m▓\033[38;5;220;48;5;94m▒\033[38;5;220;48;5;58m▒\033[38;5;178;48;5;58m░\033[38;5;178;48;5;58m░\033[38;5;136;48;5;58m░\033[38;5;221;48;5;235m░\033[38;5;222;48;5;234m \033[38;5;222;48;5;235m░\033[38;5;179;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;179;48;5;95m▒\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;173m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;130m▒\033[38;5;208;48;5;130m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;52m \033[38;5;166;48;5;234m \033[38;5;166;48;5;234m \033[38;5;130;48;5;234m \033[38;5;172;48;5;234m \033[38;5;222;48;5;235m \033[38;5;214;48;5;235m \033[38;5;214;48;5;235m \033[38;5;222;48;5;235m░\033[38;5;222;48;5;58m░\033[38;5;222;48;5;58m░\033[38;5;214;48;5;58m░\033[38;5;222;48;5;58m░\033[38;5;214;48;5;58m░\033[38;5;222;48;5;58m░\033[38;5;222;48;5;58m░\033[38;5;77;48;5;58m░\033[38;5;86;48;5;101m▒\033[38;5;167;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;236m▒\033[38;5;87;48;5;254m░\033[38;5;44;48;5;187m░\033[38;5;77;48;5;144m░\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;220;48;5;143m▓\033[38;5;220;48;5;137m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;101m▒\033[38;5;143;48;5;95m▒\033[38;5;220;48;5;240m▒\033[38;5;220;48;5;58m▒\033[38;5;220;48;5;58m▒\033[38;5;220;48;5;58m▒\033[38;5;220;48;5;94m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;220;48;5;101m▒\033[38;5;178;48;5;94m▒\033[38;5;178;48;5;58m░\033[38;5;136;48;5;58m░\033[38;5;136;48;5;58m \033[38;5;222;48;5;234m \033[38;5;172;48;5;234m \033[38;5;94;48;5;235m \033[38;5;214;48;5;58m▒\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;101m▓\033[38;5;221;48;5;101m▓\033[38;5;94;48;5;101m▓\033[38;5;214;48;5;137m▓\033[38;5;221;48;5;137m▓\033[38;5;221;48;5;101m▓\033[38;5;221;48;5;101m▓\033[38;5;94;48;5;101m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;131m▒\033[38;5;208;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;52m░\033[38;5;166;48;5;234m \033[38;5;215;48;5;234m \033[38;5;130;48;5;234m \033[38;5;172;48;5;234m \033[38;5;172;48;5;235m \033[38;5;222;48;5;235m \033[38;5;214;48;5;235m░\033[38;5;222;48;5;235m░\033[38;5;222;48;5;236m░\033[38;5;222;48;5;235m░\033[38;5;222;48;5;235m \033[38;5;94;48;5;235m \033[38;5;221;48;5;235m░\033[38;5;77;48;5;235m░\033[38;5;50;48;5;95m▒\033[38;5;209;48;5;237m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;253m░\033[38;5;178;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;144;48;5;143m▓\033[38;5;144;48;5;143m▓\033[38;5;144;48;5;137m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;95m▓\033[38;5;178;48;5;95m▓\033[38;5;178;48;5;95m▓\033[38;5;220;48;5;240m▓\033[38;5;178;48;5;240m▓\033[38;5;84;48;5;240m░\033[38;5;80;48;5;101m░\033[38;5;50;48;5;144m▒\033[38;5;50;48;5;180m▒\033[38;5;50;48;5;143m░\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;178;48;5;101m▒\033[38;5;220;48;5;58m▒\033[38;5;178;48;5;58m▒\033[38;5;136;48;5;58m░\033[38;5;136;48;5;58m░\033[38;5;221;48;5;58m▒\033[38;5;221;48;5;95m▒\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;214;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;136;48;5;137m▓\033[38;5;221;48;5;137m▓\033[38;5;221;48;5;137m▓\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;52m░\033[38;5;166;48;5;234m \033[38;5;215;48;5;234m \033[38;5;130;48;5;234m \033[38;5;172;48;5;234m \033[38;5;172;48;5;234m \033[38;5;172;48;5;235m \033[38;5;222;48;5;235m \033[38;5;222;48;5;235m░\033[38;5;214;48;5;235m░\033[38;5;222;48;5;235m░\033[38;5;130;48;5;233m \033[38;5;161;48;5;234m▓\033[38;5;43;48;5;101m▓\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;246m▒\033[38;5;220;48;5;235m▒\033[38;5;144;48;5;240m▓\033[38;5;144;48;5;101m▓\033[38;5;143;48;5;240m▒\033[38;5;185;48;5;235m░\033[38;5;185;48;5;236m▒\033[38;5;143;48;5;240m▓\033[38;5;130;48;5;241m░\033[38;5;80;48;5;101m░\033[38;5;116;48;5;144m▒\033[38;5;66;48;5;102m▓\033[38;5;174;48;5;234m▒\033[38;5;174;48;5;235m▒\033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;43;48;5;180m░\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;136;48;5;101m▒\033[38;5;178;48;5;58m▒\033[38;5;220;48;5;58m▒\033[38;5;178;48;5;58m▒\033[38;5;136;48;5;58m▒\033[38;5;136;48;5;95m▒\033[38;5;136;48;5;101m▒\033[38;5;221;48;5;101m▓\033[38;5;94;48;5;137m▓\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;214;48;5;137m▓\033[38;5;94;48;5;143m▓\033[38;5;136;48;5;143m▓\033[38;5;136;48;5;143m▓\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;58m░\033[38;5;215;48;5;234m \033[38;5;208;48;5;234m \033[38;5;130;48;5;234m \033[38;5;130;48;5;234m \033[38;5;172;48;5;234m \033[38;5;222;48;5;234m \033[38;5;222;48;5;234m \033[38;5;222;48;5;234m \033[38;5;179;48;5;235m░\033[38;5;218;48;5;238m░\033[38;5;42;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;239m▓\033[38;5;73;48;5;249m▒\033[38;5;73;48;5;246m▓\033[38;5;116;48;5;250m▒\033[38;5;73;48;5;246m▓\033[38;5;109;48;5;243m▓\033[38;5;109;48;5;244m▓\033[38;5;73;48;5;250m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m▒\033[38;5;83;48;5;137m░\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;101m▒\033[38;5;221;48;5;94m▒\033[38;5;136;48;5;58m▒\033[38;5;136;48;5;58m░\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;94m▒\033[38;5;136;48;5;101m▒\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;235m \033[38;5;215;48;5;234m \033[38;5;215;48;5;233m \033[38;5;130;48;5;233m \033[38;5;172;48;5;234m \033[38;5;172;48;5;233m \033[38;5;172;48;5;235m▒\033[38;5;103;48;5;236m▓\033[38;5;36;48;5;95m▒\033[38;5;50;48;5;145m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;86;48;5;95m▓\033[38;5;76;48;5;101m░\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;100m▒\033[38;5;221;48;5;94m▒\033[38;5;136;48;5;58m░\033[38;5;178;48;5;58m░\033[38;5;220;48;5;58m░\033[38;5;178;48;5;94m▒\033[38;5;178;48;5;101m▒\033[38;5;136;48;5;137m▓\033[38;5;136;48;5;143m▓\033[38;5;221;48;5;143m▓\033[38;5;94;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;179;48;5;144m▒\033[38;5;172;48;5;144m▒\033[38;5;172;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;221;48;5;143m▓\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;234m \033[38;5;166;48;5;233m \033[38;5;215;48;5;233m \033[38;5;166;48;5;233m \033[38;5;130;48;5;233m \033[38;5;112;48;5;236m░\033[38;5;43;48;5;59m▓\033[38;5;84;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;235m▒\033[38;5;79;48;5;243m▓\033[38;5;73;48;5;144m▒\033[38;5;80;48;5;144m▒\033[38;5;31;48;5;101m▓\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;136m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;94m▒\033[38;5;221;48;5;58m▒\033[38;5;136;48;5;58m▒\033[38;5;178;48;5;101m▒\033[38;5;136;48;5;137m▓\033[38;5;221;48;5;144m▓\033[38;5;221;48;5;144m▒\033[38;5;94;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;221;48;5;137m▓\033[38;5;136;48;5;137m▓\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;130;48;5;236m░\033[38;5;166;48;5;233m \033[38;5;166;48;5;233m \033[38;5;174;48;5;237m▒\033[38;5;220;48;5;238m▓\033[38;5;174;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;249m▒\033[38;5;116;48;5;144m▒\033[38;5;80;48;5;181m░\033[38;5;153;48;5;144m░\033[38;5;81;48;5;101m░\033[38;5;94;48;5;101m▓\033[38;5;214;48;5;95m▓\033[38;5;179;48;5;95m▒\033[38;5;94;48;5;94m▒\033[38;5;221;48;5;3m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;136;48;5;101m▒\033[38;5;50;48;5;137m░\033[38;5;50;48;5;137m▒\033[38;5;50;48;5;101m░\033[38;5;29;48;5;95m▓\033[38;5;32;48;5;101m▒\033[38;5;27;48;5;138m▒\033[38;5;57;48;5;144m░\033[38;5;94;48;5;181m▓\033[38;5;136;48;5;181m▓\033[38;5;94;48;5;181m▓\033[38;5;94;48;5;181m▓\033[38;5;94;48;5;181m▓\033[38;5;179;48;5;180m▓\033[38;5;221;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;221;48;5;144m▓\033[38;5;136;48;5;144m▓\033[38;5;178;48;5;144m▓\033[38;5;136;48;5;137m▓\033[38;5;178;48;5;101m▓\033[38;5;178;48;5;95m▓\033[38;5;221;48;5;58m▒\033[38;5;94;48;5;101m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;180;48;5;58m▒\033[38;5;180;48;5;237m▒\033[38;5;137;48;5;237m▒\033[38;5;50;48;5;241m▒\033[38;5;50;48;5;248m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;171;48;5;101m░\033[38;5;119;48;5;101m░\033[38;5;178;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;101m▒\033[38;5;136;48;5;101m▒\033[38;5;136;48;5;101m▒\033[38;5;221;48;5;95m▒\033[38;5;221;48;5;95m▒\033[38;5;136;48;5;101m▒\033[38;5;178;48;5;137m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;178;48;5;137m▓\033[38;5;50;48;5;144m▒\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;116;48;5;187m▒\033[38;5;73;48;5;144m▒\033[38;5;50;48;5;137m▒\033[38;5;110;48;5;95m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;180;48;5;58m▒\033[38;5;208;48;5;236m▒\033[38;5;43;48;5;240m░\033[38;5;209;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;246m▓\033[38;5;21;48;5;238m░\033[38;5;220;48;5;233m \033[38;5;220;48;5;235m░\033[38;5;136;48;5;58m▒\033[38;5;136;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;112;48;5;143m▒\033[38;5;73;48;5;246m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;236m▒\033[38;5;50;48;5;180m░\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;180;48;5;58m▒\033[38;5;43;48;5;95m░\033[38;5;86;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;246m▓\033[38;5;93;48;5;101m░\033[38;5;136;48;5;101m▓\033[38;5;178;48;5;101m▓\033[38;5;178;48;5;137m▓\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;220;48;5;179m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;86;48;5;143m░\033[38;5;80;48;5;186m▒\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;236m▒\033[38;5;50;48;5;180m░\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;38;48;5;239m▓\033[38;5;36;48;5;138m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;7m▒\033[38;5;45;48;5;95m░\033[38;5;136;48;5;101m▓\033[38;5;178;48;5;137m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▓\033[38;5;80;48;5;187m░\033[38;5;131;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;236m▒\033[38;5;50;48;5;187m░\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;36;48;5;95m░\033[38;5;50;48;5;249m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m▒\033[38;5;44;48;5;187m░\033[38;5;220;48;5;137m▓\033[38;5;220;48;5;137m▓\033[38;5;220;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;201;48;5;144m░\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;104;48;5;180m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m▒\033[38;5;200;48;5;95m▒\033[38;5;50;48;5;248m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;238m▓\033[38;5;80;48;5;144m▒\033[38;5;84;48;5;101m░\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;137m▓\033[38;5;220;48;5;101m▓\033[38;5;178;48;5;95m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;95m▒\033[38;5;220;48;5;101m▓\033[38;5;33;48;5;101m▒\033[38;5;50;48;5;137m░\033[38;5;50;48;5;181m▒\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;117;48;5;144m░\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;180;48;5;58m▒\033[38;5;119;48;5;95m░\033[38;5;50;48;5;247m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;204;48;5;236m▒\033[38;5;204;48;5;237m▒\033[38;5;204;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;224m░\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;220;48;5;95m▒\033[38;5;50;48;5;247m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;246m▓\033[38;5;50;48;5;181m░\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;172;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;43;48;5;101m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;245m▓\033[38;5;84;48;5;180m░\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;58m░\033[38;5;119;48;5;239m░\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m░\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;94;48;5;95m░\033[38;5;209;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[38;5;80;48;5;187m░\033[38;5;136;48;5;144m▓\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;43;48;5;138m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m▒\033[38;5;136;48;5;144m▓\033[38;5;214;48;5;137m▓\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;179m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m░\033[38;5;19;48;5;94m░\033[38;5;50;48;5;181m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;236m▒\033[38;5;80;48;5;246m░\033[38;5;179;48;5;101m▓\033[38;5;172;48;5;137m▓\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;95m▒\033[38;5;214;48;5;95m▒\033[38;5;50;48;5;101m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;244m▒\033[38;5;214;48;5;238m▓\033[38;5;179;48;5;95m▓\033[38;5;94;48;5;240m▒\033[38;5;94;48;5;95m▓\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;95m▓\033[38;5;34;48;5;237m░\033[38;5;80;48;5;59m░\033[38;5;116;48;5;250m▒\033[38;5;138;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
        $display("\033[0m");
    endtask

    initial begin
        i_rst_n = 1'b1;
        i_start = 1'b0;
        i_pause = 1'b0;
        i_speed = `SPEED - 1;
        i_is_slow = `IS_SLOW;
        i_slow_mode = `SLOW_MODE;
        i_daclrck = 1'b0;
        i_sram_data = 16'h0000;
        i_sram_stop_addr = 20'hfffff;

        error = 0;
        diff = 0;
        
        // 加載記憶體數據
        load_mem_data(`MEMFILE, fp_mem, mem_data);
        
        // 加載 golden 數據
        load_golden_data(`GOLDENFILE, fp_golden, golden_data);

        // Reset sequence
        #(`CYCLE * 2.5) i_rst_n = 1'b0;
        #(`CYCLE * 3) i_rst_n = 1'b1;
        #(`CYCLE * 1) i_start = 1'b1;
        #(`CYCLE * 2) i_start = 1'b0;
        #(`CYCLE * 2) i_pause = 1'b1;
        #(`CYCLE * 1) i_pause = 1'b0;

        @(posedge i_clk) i_daclrck = 1'b1;
        // repeat (100) begin
        //     #(`CYCLE * 20) i_daclrck = 1'b0;
        //     #(`CYCLE * 20) i_daclrck = 1'b1;
        // end
        for (i = 0; i < `SIM_CYCLES; i = i + 1) begin
            i_sram_data = mem_data[o_sram_addr];
            #(`CYCLE * 20);
            i_daclrck = 1'b0;
            diff = o_dac_data - golden_data[i];
            if(o_en) begin
                if(diff < -1 || diff > 1) begin
                    // ignore diff = 1 or -1, we can accept this error
                    $display("Diff bigger than 1: Mismatch at case %d", i);
                    $display("Golden: %16b", golden_data[i]);
                    $display("Output: %16b", o_dac_data);
                    $display("");
                    error = error + 1;
                end
            end
            #(`CYCLE * 20);
            i_daclrck = 1'b1;
        end

        if (error == 0) begin
            display_graph_pass;
            $display("==========================================");
            $display("======  Congratulations! You Pass!  ======");
            $display("==========================================");
        end else begin
            display_graph_fail;
            $display("===============================");
            $display("There are %0d errors.", error);
            $display("===============================");
        end
        

        $finish;
    end

    initial begin
        $fsdbDumpfile("tb_AudDSP.fsdb");
        $fsdbDumpvars;
    end
    // initial #(`CYCLE*10000000) $finish;
endmodule