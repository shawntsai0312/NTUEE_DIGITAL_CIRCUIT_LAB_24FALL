module SramDecoder (
    input i_clk,
    input i_rst_n,
    input [11:0] VGA_H_pos,
    input [11:0] VGA_V_pos,
    input [11:0] Car_x,
    input [11:0] Car_y,
    output [23:0] o_color
);

endmodule