module image_data(output reg [2:0] pixel_data [0:1599]);
    initial begin
        pixel_data[0] = 3'b011; // x=0, y=0
        pixel_data[1] = 3'b010; // x=1, y=0
        pixel_data[2] = 3'b010; // x=2, y=0
        pixel_data[3] = 3'b010; // x=3, y=0
        pixel_data[4] = 3'b010; // x=4, y=0
        pixel_data[5] = 3'b010; // x=5, y=0
        pixel_data[6] = 3'b010; // x=6, y=0
        pixel_data[7] = 3'b010; // x=7, y=0
        pixel_data[8] = 3'b010; // x=8, y=0
        pixel_data[9] = 3'b011; // x=9, y=0
        pixel_data[10] = 3'b010; // x=10, y=0
        pixel_data[11] = 3'b010; // x=11, y=0
        pixel_data[12] = 3'b010; // x=12, y=0
        pixel_data[13] = 3'b010; // x=13, y=0
        pixel_data[14] = 3'b010; // x=14, y=0
        pixel_data[15] = 3'b010; // x=15, y=0
        pixel_data[16] = 3'b010; // x=16, y=0
        pixel_data[17] = 3'b010; // x=17, y=0
        pixel_data[18] = 3'b010; // x=18, y=0
        pixel_data[19] = 3'b010; // x=19, y=0
        pixel_data[20] = 3'b011; // x=20, y=0
        pixel_data[21] = 3'b010; // x=21, y=0
        pixel_data[22] = 3'b010; // x=22, y=0
        pixel_data[23] = 3'b010; // x=23, y=0
        pixel_data[24] = 3'b010; // x=24, y=0
        pixel_data[25] = 3'b010; // x=25, y=0
        pixel_data[26] = 3'b010; // x=26, y=0
        pixel_data[27] = 3'b010; // x=27, y=0
        pixel_data[28] = 3'b010; // x=28, y=0
        pixel_data[29] = 3'b010; // x=29, y=0
        pixel_data[30] = 3'b010; // x=30, y=0
        pixel_data[31] = 3'b010; // x=31, y=0
        pixel_data[32] = 3'b010; // x=32, y=0
        pixel_data[33] = 3'b011; // x=33, y=0
        pixel_data[34] = 3'b010; // x=34, y=0
        pixel_data[35] = 3'b010; // x=35, y=0
        pixel_data[36] = 3'b010; // x=36, y=0
        pixel_data[37] = 3'b010; // x=37, y=0
        pixel_data[38] = 3'b010; // x=38, y=0
        pixel_data[39] = 3'b010; // x=39, y=0
        pixel_data[40] = 3'b010; // x=0, y=1
        pixel_data[41] = 3'b011; // x=1, y=1
        pixel_data[42] = 3'b010; // x=2, y=1
        pixel_data[43] = 3'b010; // x=3, y=1
        pixel_data[44] = 3'b010; // x=4, y=1
        pixel_data[45] = 3'b010; // x=5, y=1
        pixel_data[46] = 3'b010; // x=6, y=1
        pixel_data[47] = 3'b010; // x=7, y=1
        pixel_data[48] = 3'b010; // x=8, y=1
        pixel_data[49] = 3'b010; // x=9, y=1
        pixel_data[50] = 3'b010; // x=10, y=1
        pixel_data[51] = 3'b010; // x=11, y=1
        pixel_data[52] = 3'b010; // x=12, y=1
        pixel_data[53] = 3'b010; // x=13, y=1
        pixel_data[54] = 3'b010; // x=14, y=1
        pixel_data[55] = 3'b010; // x=15, y=1
        pixel_data[56] = 3'b010; // x=16, y=1
        pixel_data[57] = 3'b010; // x=17, y=1
        pixel_data[58] = 3'b010; // x=18, y=1
        pixel_data[59] = 3'b011; // x=19, y=1
        pixel_data[60] = 3'b010; // x=20, y=1
        pixel_data[61] = 3'b010; // x=21, y=1
        pixel_data[62] = 3'b010; // x=22, y=1
        pixel_data[63] = 3'b011; // x=23, y=1
        pixel_data[64] = 3'b010; // x=24, y=1
        pixel_data[65] = 3'b010; // x=25, y=1
        pixel_data[66] = 3'b010; // x=26, y=1
        pixel_data[67] = 3'b010; // x=27, y=1
        pixel_data[68] = 3'b010; // x=28, y=1
        pixel_data[69] = 3'b010; // x=29, y=1
        pixel_data[70] = 3'b011; // x=30, y=1
        pixel_data[71] = 3'b010; // x=31, y=1
        pixel_data[72] = 3'b010; // x=32, y=1
        pixel_data[73] = 3'b010; // x=33, y=1
        pixel_data[74] = 3'b011; // x=34, y=1
        pixel_data[75] = 3'b010; // x=35, y=1
        pixel_data[76] = 3'b010; // x=36, y=1
        pixel_data[77] = 3'b010; // x=37, y=1
        pixel_data[78] = 3'b010; // x=38, y=1
        pixel_data[79] = 3'b010; // x=39, y=1
        pixel_data[80] = 3'b010; // x=0, y=2
        pixel_data[81] = 3'b010; // x=1, y=2
        pixel_data[82] = 3'b011; // x=2, y=2
        pixel_data[83] = 3'b010; // x=3, y=2
        pixel_data[84] = 3'b010; // x=4, y=2
        pixel_data[85] = 3'b010; // x=5, y=2
        pixel_data[86] = 3'b010; // x=6, y=2
        pixel_data[87] = 3'b010; // x=7, y=2
        pixel_data[88] = 3'b011; // x=8, y=2
        pixel_data[89] = 3'b010; // x=9, y=2
        pixel_data[90] = 3'b010; // x=10, y=2
        pixel_data[91] = 3'b010; // x=11, y=2
        pixel_data[92] = 3'b010; // x=12, y=2
        pixel_data[93] = 3'b011; // x=13, y=2
        pixel_data[94] = 3'b010; // x=14, y=2
        pixel_data[95] = 3'b010; // x=15, y=2
        pixel_data[96] = 3'b010; // x=16, y=2
        pixel_data[97] = 3'b010; // x=17, y=2
        pixel_data[98] = 3'b010; // x=18, y=2
        pixel_data[99] = 3'b010; // x=19, y=2
        pixel_data[100] = 3'b010; // x=20, y=2
        pixel_data[101] = 3'b010; // x=21, y=2
        pixel_data[102] = 3'b010; // x=22, y=2
        pixel_data[103] = 3'b010; // x=23, y=2
        pixel_data[104] = 3'b011; // x=24, y=2
        pixel_data[105] = 3'b010; // x=25, y=2
        pixel_data[106] = 3'b010; // x=26, y=2
        pixel_data[107] = 3'b010; // x=27, y=2
        pixel_data[108] = 3'b010; // x=28, y=2
        pixel_data[109] = 3'b010; // x=29, y=2
        pixel_data[110] = 3'b010; // x=30, y=2
        pixel_data[111] = 3'b010; // x=31, y=2
        pixel_data[112] = 3'b010; // x=32, y=2
        pixel_data[113] = 3'b010; // x=33, y=2
        pixel_data[114] = 3'b010; // x=34, y=2
        pixel_data[115] = 3'b010; // x=35, y=2
        pixel_data[116] = 3'b010; // x=36, y=2
        pixel_data[117] = 3'b010; // x=37, y=2
        pixel_data[118] = 3'b010; // x=38, y=2
        pixel_data[119] = 3'b010; // x=39, y=2
        pixel_data[120] = 3'b010; // x=0, y=3
        pixel_data[121] = 3'b010; // x=1, y=3
        pixel_data[122] = 3'b010; // x=2, y=3
        pixel_data[123] = 3'b011; // x=3, y=3
        pixel_data[124] = 3'b010; // x=4, y=3
        pixel_data[125] = 3'b010; // x=5, y=3
        pixel_data[126] = 3'b011; // x=6, y=3
        pixel_data[127] = 3'b011; // x=7, y=3
        pixel_data[128] = 3'b010; // x=8, y=3
        pixel_data[129] = 3'b010; // x=9, y=3
        pixel_data[130] = 3'b010; // x=10, y=3
        pixel_data[131] = 3'b010; // x=11, y=3
        pixel_data[132] = 3'b010; // x=12, y=3
        pixel_data[133] = 3'b010; // x=13, y=3
        pixel_data[134] = 3'b011; // x=14, y=3
        pixel_data[135] = 3'b010; // x=15, y=3
        pixel_data[136] = 3'b010; // x=16, y=3
        pixel_data[137] = 3'b011; // x=17, y=3
        pixel_data[138] = 3'b010; // x=18, y=3
        pixel_data[139] = 3'b010; // x=19, y=3
        pixel_data[140] = 3'b010; // x=20, y=3
        pixel_data[141] = 3'b010; // x=21, y=3
        pixel_data[142] = 3'b010; // x=22, y=3
        pixel_data[143] = 3'b010; // x=23, y=3
        pixel_data[144] = 3'b010; // x=24, y=3
        pixel_data[145] = 3'b011; // x=25, y=3
        pixel_data[146] = 3'b010; // x=26, y=3
        pixel_data[147] = 3'b011; // x=27, y=3
        pixel_data[148] = 3'b011; // x=28, y=3
        pixel_data[149] = 3'b010; // x=29, y=3
        pixel_data[150] = 3'b010; // x=30, y=3
        pixel_data[151] = 3'b010; // x=31, y=3
        pixel_data[152] = 3'b010; // x=32, y=3
        pixel_data[153] = 3'b010; // x=33, y=3
        pixel_data[154] = 3'b010; // x=34, y=3
        pixel_data[155] = 3'b010; // x=35, y=3
        pixel_data[156] = 3'b011; // x=36, y=3
        pixel_data[157] = 3'b010; // x=37, y=3
        pixel_data[158] = 3'b011; // x=38, y=3
        pixel_data[159] = 3'b011; // x=39, y=3
        pixel_data[160] = 3'b010; // x=0, y=4
        pixel_data[161] = 3'b010; // x=1, y=4
        pixel_data[162] = 3'b010; // x=2, y=4
        pixel_data[163] = 3'b010; // x=3, y=4
        pixel_data[164] = 3'b010; // x=4, y=4
        pixel_data[165] = 3'b011; // x=5, y=4
        pixel_data[166] = 3'b011; // x=6, y=4
        pixel_data[167] = 3'b010; // x=7, y=4
        pixel_data[168] = 3'b010; // x=8, y=4
        pixel_data[169] = 3'b010; // x=9, y=4
        pixel_data[170] = 3'b010; // x=10, y=4
        pixel_data[171] = 3'b010; // x=11, y=4
        pixel_data[172] = 3'b010; // x=12, y=4
        pixel_data[173] = 3'b010; // x=13, y=4
        pixel_data[174] = 3'b010; // x=14, y=4
        pixel_data[175] = 3'b010; // x=15, y=4
        pixel_data[176] = 3'b011; // x=16, y=4
        pixel_data[177] = 3'b011; // x=17, y=4
        pixel_data[178] = 3'b010; // x=18, y=4
        pixel_data[179] = 3'b010; // x=19, y=4
        pixel_data[180] = 3'b010; // x=20, y=4
        pixel_data[181] = 3'b010; // x=21, y=4
        pixel_data[182] = 3'b010; // x=22, y=4
        pixel_data[183] = 3'b010; // x=23, y=4
        pixel_data[184] = 3'b010; // x=24, y=4
        pixel_data[185] = 3'b010; // x=25, y=4
        pixel_data[186] = 3'b011; // x=26, y=4
        pixel_data[187] = 3'b011; // x=27, y=4
        pixel_data[188] = 3'b011; // x=28, y=4
        pixel_data[189] = 3'b010; // x=29, y=4
        pixel_data[190] = 3'b010; // x=30, y=4
        pixel_data[191] = 3'b010; // x=31, y=4
        pixel_data[192] = 3'b010; // x=32, y=4
        pixel_data[193] = 3'b010; // x=33, y=4
        pixel_data[194] = 3'b010; // x=34, y=4
        pixel_data[195] = 3'b010; // x=35, y=4
        pixel_data[196] = 3'b010; // x=36, y=4
        pixel_data[197] = 3'b011; // x=37, y=4
        pixel_data[198] = 3'b011; // x=38, y=4
        pixel_data[199] = 3'b011; // x=39, y=4
        pixel_data[200] = 3'b010; // x=0, y=5
        pixel_data[201] = 3'b010; // x=1, y=5
        pixel_data[202] = 3'b010; // x=2, y=5
        pixel_data[203] = 3'b010; // x=3, y=5
        pixel_data[204] = 3'b011; // x=4, y=5
        pixel_data[205] = 3'b011; // x=5, y=5
        pixel_data[206] = 3'b011; // x=6, y=5
        pixel_data[207] = 3'b010; // x=7, y=5
        pixel_data[208] = 3'b010; // x=8, y=5
        pixel_data[209] = 3'b010; // x=9, y=5
        pixel_data[210] = 3'b010; // x=10, y=5
        pixel_data[211] = 3'b010; // x=11, y=5
        pixel_data[212] = 3'b010; // x=12, y=5
        pixel_data[213] = 3'b010; // x=13, y=5
        pixel_data[214] = 3'b010; // x=14, y=5
        pixel_data[215] = 3'b011; // x=15, y=5
        pixel_data[216] = 3'b011; // x=16, y=5
        pixel_data[217] = 3'b011; // x=17, y=5
        pixel_data[218] = 3'b010; // x=18, y=5
        pixel_data[219] = 3'b010; // x=19, y=5
        pixel_data[220] = 3'b010; // x=20, y=5
        pixel_data[221] = 3'b010; // x=21, y=5
        pixel_data[222] = 3'b010; // x=22, y=5
        pixel_data[223] = 3'b010; // x=23, y=5
        pixel_data[224] = 3'b010; // x=24, y=5
        pixel_data[225] = 3'b010; // x=25, y=5
        pixel_data[226] = 3'b011; // x=26, y=5
        pixel_data[227] = 3'b011; // x=27, y=5
        pixel_data[228] = 3'b011; // x=28, y=5
        pixel_data[229] = 3'b010; // x=29, y=5
        pixel_data[230] = 3'b010; // x=30, y=5
        pixel_data[231] = 3'b010; // x=31, y=5
        pixel_data[232] = 3'b010; // x=32, y=5
        pixel_data[233] = 3'b010; // x=33, y=5
        pixel_data[234] = 3'b010; // x=34, y=5
        pixel_data[235] = 3'b010; // x=35, y=5
        pixel_data[236] = 3'b011; // x=36, y=5
        pixel_data[237] = 3'b011; // x=37, y=5
        pixel_data[238] = 3'b011; // x=38, y=5
        pixel_data[239] = 3'b010; // x=39, y=5
        pixel_data[240] = 3'b010; // x=0, y=6
        pixel_data[241] = 3'b010; // x=1, y=6
        pixel_data[242] = 3'b001; // x=2, y=6
        pixel_data[243] = 3'b011; // x=3, y=6
        pixel_data[244] = 3'b011; // x=4, y=6
        pixel_data[245] = 3'b011; // x=5, y=6
        pixel_data[246] = 3'b010; // x=6, y=6
        pixel_data[247] = 3'b010; // x=7, y=6
        pixel_data[248] = 3'b010; // x=8, y=6
        pixel_data[249] = 3'b010; // x=9, y=6
        pixel_data[250] = 3'b010; // x=10, y=6
        pixel_data[251] = 3'b010; // x=11, y=6
        pixel_data[252] = 3'b010; // x=12, y=6
        pixel_data[253] = 3'b010; // x=13, y=6
        pixel_data[254] = 3'b011; // x=14, y=6
        pixel_data[255] = 3'b011; // x=15, y=6
        pixel_data[256] = 3'b011; // x=16, y=6
        pixel_data[257] = 3'b010; // x=17, y=6
        pixel_data[258] = 3'b010; // x=18, y=6
        pixel_data[259] = 3'b010; // x=19, y=6
        pixel_data[260] = 3'b010; // x=20, y=6
        pixel_data[261] = 3'b010; // x=21, y=6
        pixel_data[262] = 3'b010; // x=22, y=6
        pixel_data[263] = 3'b010; // x=23, y=6
        pixel_data[264] = 3'b010; // x=24, y=6
        pixel_data[265] = 3'b011; // x=25, y=6
        pixel_data[266] = 3'b011; // x=26, y=6
        pixel_data[267] = 3'b011; // x=27, y=6
        pixel_data[268] = 3'b010; // x=28, y=6
        pixel_data[269] = 3'b010; // x=29, y=6
        pixel_data[270] = 3'b010; // x=30, y=6
        pixel_data[271] = 3'b010; // x=31, y=6
        pixel_data[272] = 3'b010; // x=32, y=6
        pixel_data[273] = 3'b010; // x=33, y=6
        pixel_data[274] = 3'b010; // x=34, y=6
        pixel_data[275] = 3'b010; // x=35, y=6
        pixel_data[276] = 3'b011; // x=36, y=6
        pixel_data[277] = 3'b011; // x=37, y=6
        pixel_data[278] = 3'b011; // x=38, y=6
        pixel_data[279] = 3'b010; // x=39, y=6
        pixel_data[280] = 3'b010; // x=0, y=7
        pixel_data[281] = 3'b010; // x=1, y=7
        pixel_data[282] = 3'b010; // x=2, y=7
        pixel_data[283] = 3'b011; // x=3, y=7
        pixel_data[284] = 3'b010; // x=4, y=7
        pixel_data[285] = 3'b010; // x=5, y=7
        pixel_data[286] = 3'b010; // x=6, y=7
        pixel_data[287] = 3'b011; // x=7, y=7
        pixel_data[288] = 3'b010; // x=8, y=7
        pixel_data[289] = 3'b010; // x=9, y=7
        pixel_data[290] = 3'b010; // x=10, y=7
        pixel_data[291] = 3'b010; // x=11, y=7
        pixel_data[292] = 3'b010; // x=12, y=7
        pixel_data[293] = 3'b010; // x=13, y=7
        pixel_data[294] = 3'b011; // x=14, y=7
        pixel_data[295] = 3'b010; // x=15, y=7
        pixel_data[296] = 3'b010; // x=16, y=7
        pixel_data[297] = 3'b010; // x=17, y=7
        pixel_data[298] = 3'b011; // x=18, y=7
        pixel_data[299] = 3'b010; // x=19, y=7
        pixel_data[300] = 3'b010; // x=20, y=7
        pixel_data[301] = 3'b010; // x=21, y=7
        pixel_data[302] = 3'b010; // x=22, y=7
        pixel_data[303] = 3'b010; // x=23, y=7
        pixel_data[304] = 3'b010; // x=24, y=7
        pixel_data[305] = 3'b011; // x=25, y=7
        pixel_data[306] = 3'b010; // x=26, y=7
        pixel_data[307] = 3'b010; // x=27, y=7
        pixel_data[308] = 3'b010; // x=28, y=7
        pixel_data[309] = 3'b011; // x=29, y=7
        pixel_data[310] = 3'b010; // x=30, y=7
        pixel_data[311] = 3'b010; // x=31, y=7
        pixel_data[312] = 3'b010; // x=32, y=7
        pixel_data[313] = 3'b010; // x=33, y=7
        pixel_data[314] = 3'b010; // x=34, y=7
        pixel_data[315] = 3'b010; // x=35, y=7
        pixel_data[316] = 3'b011; // x=36, y=7
        pixel_data[317] = 3'b010; // x=37, y=7
        pixel_data[318] = 3'b010; // x=38, y=7
        pixel_data[319] = 3'b010; // x=39, y=7
        pixel_data[320] = 3'b010; // x=0, y=8
        pixel_data[321] = 3'b010; // x=1, y=8
        pixel_data[322] = 3'b011; // x=2, y=8
        pixel_data[323] = 3'b010; // x=3, y=8
        pixel_data[324] = 3'b010; // x=4, y=8
        pixel_data[325] = 3'b010; // x=5, y=8
        pixel_data[326] = 3'b010; // x=6, y=8
        pixel_data[327] = 3'b010; // x=7, y=8
        pixel_data[328] = 3'b011; // x=8, y=8
        pixel_data[329] = 3'b010; // x=9, y=8
        pixel_data[330] = 3'b010; // x=10, y=8
        pixel_data[331] = 3'b010; // x=11, y=8
        pixel_data[332] = 3'b010; // x=12, y=8
        pixel_data[333] = 3'b010; // x=13, y=8
        pixel_data[334] = 3'b010; // x=14, y=8
        pixel_data[335] = 3'b001; // x=15, y=8
        pixel_data[336] = 3'b000; // x=16, y=8
        pixel_data[337] = 3'b010; // x=17, y=8
        pixel_data[338] = 3'b010; // x=18, y=8
        pixel_data[339] = 3'b011; // x=19, y=8
        pixel_data[340] = 3'b010; // x=20, y=8
        pixel_data[341] = 3'b010; // x=21, y=8
        pixel_data[342] = 3'b010; // x=22, y=8
        pixel_data[343] = 3'b010; // x=23, y=8
        pixel_data[344] = 3'b010; // x=24, y=8
        pixel_data[345] = 3'b010; // x=25, y=8
        pixel_data[346] = 3'b010; // x=26, y=8
        pixel_data[347] = 3'b010; // x=27, y=8
        pixel_data[348] = 3'b010; // x=28, y=8
        pixel_data[349] = 3'b010; // x=29, y=8
        pixel_data[350] = 3'b011; // x=30, y=8
        pixel_data[351] = 3'b010; // x=31, y=8
        pixel_data[352] = 3'b010; // x=32, y=8
        pixel_data[353] = 3'b010; // x=33, y=8
        pixel_data[354] = 3'b011; // x=34, y=8
        pixel_data[355] = 3'b011; // x=35, y=8
        pixel_data[356] = 3'b010; // x=36, y=8
        pixel_data[357] = 3'b010; // x=37, y=8
        pixel_data[358] = 3'b010; // x=38, y=8
        pixel_data[359] = 3'b010; // x=39, y=8
        pixel_data[360] = 3'b010; // x=0, y=9
        pixel_data[361] = 3'b011; // x=1, y=9
        pixel_data[362] = 3'b010; // x=2, y=9
        pixel_data[363] = 3'b010; // x=3, y=9
        pixel_data[364] = 3'b010; // x=4, y=9
        pixel_data[365] = 3'b010; // x=5, y=9
        pixel_data[366] = 3'b010; // x=6, y=9
        pixel_data[367] = 3'b001; // x=7, y=9
        pixel_data[368] = 3'b010; // x=8, y=9
        pixel_data[369] = 3'b010; // x=9, y=9
        pixel_data[370] = 3'b001; // x=10, y=9
        pixel_data[371] = 3'b010; // x=11, y=9
        pixel_data[372] = 3'b010; // x=12, y=9
        pixel_data[373] = 3'b001; // x=13, y=9
        pixel_data[374] = 3'b000; // x=14, y=9
        pixel_data[375] = 3'b100; // x=15, y=9
        pixel_data[376] = 3'b100; // x=16, y=9
        pixel_data[377] = 3'b000; // x=17, y=9
        pixel_data[378] = 3'b001; // x=18, y=9
        pixel_data[379] = 3'b001; // x=19, y=9
        pixel_data[380] = 3'b001; // x=20, y=9
        pixel_data[381] = 3'b001; // x=21, y=9
        pixel_data[382] = 3'b000; // x=22, y=9
        pixel_data[383] = 3'b000; // x=23, y=9
        pixel_data[384] = 3'b001; // x=24, y=9
        pixel_data[385] = 3'b000; // x=25, y=9
        pixel_data[386] = 3'b000; // x=26, y=9
        pixel_data[387] = 3'b001; // x=27, y=9
        pixel_data[388] = 3'b001; // x=28, y=9
        pixel_data[389] = 3'b010; // x=29, y=9
        pixel_data[390] = 3'b010; // x=30, y=9
        pixel_data[391] = 3'b010; // x=31, y=9
        pixel_data[392] = 3'b010; // x=32, y=9
        pixel_data[393] = 3'b010; // x=33, y=9
        pixel_data[394] = 3'b010; // x=34, y=9
        pixel_data[395] = 3'b010; // x=35, y=9
        pixel_data[396] = 3'b010; // x=36, y=9
        pixel_data[397] = 3'b010; // x=37, y=9
        pixel_data[398] = 3'b010; // x=38, y=9
        pixel_data[399] = 3'b010; // x=39, y=9
        pixel_data[400] = 3'b010; // x=0, y=10
        pixel_data[401] = 3'b010; // x=1, y=10
        pixel_data[402] = 3'b010; // x=2, y=10
        pixel_data[403] = 3'b001; // x=3, y=10
        pixel_data[404] = 3'b000; // x=4, y=10
        pixel_data[405] = 3'b000; // x=5, y=10
        pixel_data[406] = 3'b011; // x=6, y=10
        pixel_data[407] = 3'b011; // x=7, y=10
        pixel_data[408] = 3'b011; // x=8, y=10
        pixel_data[409] = 3'b011; // x=9, y=10
        pixel_data[410] = 3'b011; // x=10, y=10
        pixel_data[411] = 3'b011; // x=11, y=10
        pixel_data[412] = 3'b011; // x=12, y=10
        pixel_data[413] = 3'b011; // x=13, y=10
        pixel_data[414] = 3'b011; // x=14, y=10
        pixel_data[415] = 3'b100; // x=15, y=10
        pixel_data[416] = 3'b101; // x=16, y=10
        pixel_data[417] = 3'b000; // x=17, y=10
        pixel_data[418] = 3'b011; // x=18, y=10
        pixel_data[419] = 3'b011; // x=19, y=10
        pixel_data[420] = 3'b011; // x=20, y=10
        pixel_data[421] = 3'b011; // x=21, y=10
        pixel_data[422] = 3'b100; // x=22, y=10
        pixel_data[423] = 3'b100; // x=23, y=10
        pixel_data[424] = 3'b011; // x=24, y=10
        pixel_data[425] = 3'b100; // x=25, y=10
        pixel_data[426] = 3'b100; // x=26, y=10
        pixel_data[427] = 3'b001; // x=27, y=10
        pixel_data[428] = 3'b010; // x=28, y=10
        pixel_data[429] = 3'b000; // x=29, y=10
        pixel_data[430] = 3'b000; // x=30, y=10
        pixel_data[431] = 3'b001; // x=31, y=10
        pixel_data[432] = 3'b000; // x=32, y=10
        pixel_data[433] = 3'b000; // x=33, y=10
        pixel_data[434] = 3'b000; // x=34, y=10
        pixel_data[435] = 3'b000; // x=35, y=10
        pixel_data[436] = 3'b010; // x=36, y=10
        pixel_data[437] = 3'b010; // x=37, y=10
        pixel_data[438] = 3'b010; // x=38, y=10
        pixel_data[439] = 3'b010; // x=39, y=10
        pixel_data[440] = 3'b010; // x=0, y=11
        pixel_data[441] = 3'b010; // x=1, y=11
        pixel_data[442] = 3'b000; // x=2, y=11
        pixel_data[443] = 3'b011; // x=3, y=11
        pixel_data[444] = 3'b100; // x=4, y=11
        pixel_data[445] = 3'b101; // x=5, y=11
        pixel_data[446] = 3'b101; // x=6, y=11
        pixel_data[447] = 3'b101; // x=7, y=11
        pixel_data[448] = 3'b101; // x=8, y=11
        pixel_data[449] = 3'b101; // x=9, y=11
        pixel_data[450] = 3'b101; // x=10, y=11
        pixel_data[451] = 3'b101; // x=11, y=11
        pixel_data[452] = 3'b101; // x=12, y=11
        pixel_data[453] = 3'b101; // x=13, y=11
        pixel_data[454] = 3'b101; // x=14, y=11
        pixel_data[455] = 3'b110; // x=15, y=11
        pixel_data[456] = 3'b110; // x=16, y=11
        pixel_data[457] = 3'b110; // x=17, y=11
        pixel_data[458] = 3'b110; // x=18, y=11
        pixel_data[459] = 3'b110; // x=19, y=11
        pixel_data[460] = 3'b110; // x=20, y=11
        pixel_data[461] = 3'b110; // x=21, y=11
        pixel_data[462] = 3'b110; // x=22, y=11
        pixel_data[463] = 3'b111; // x=23, y=11
        pixel_data[464] = 3'b110; // x=24, y=11
        pixel_data[465] = 3'b110; // x=25, y=11
        pixel_data[466] = 3'b111; // x=26, y=11
        pixel_data[467] = 3'b110; // x=27, y=11
        pixel_data[468] = 3'b110; // x=28, y=11
        pixel_data[469] = 3'b110; // x=29, y=11
        pixel_data[470] = 3'b110; // x=30, y=11
        pixel_data[471] = 3'b101; // x=31, y=11
        pixel_data[472] = 3'b101; // x=32, y=11
        pixel_data[473] = 3'b101; // x=33, y=11
        pixel_data[474] = 3'b100; // x=34, y=11
        pixel_data[475] = 3'b100; // x=35, y=11
        pixel_data[476] = 3'b010; // x=36, y=11
        pixel_data[477] = 3'b001; // x=37, y=11
        pixel_data[478] = 3'b010; // x=38, y=11
        pixel_data[479] = 3'b010; // x=39, y=11
        pixel_data[480] = 3'b010; // x=0, y=12
        pixel_data[481] = 3'b001; // x=1, y=12
        pixel_data[482] = 3'b011; // x=2, y=12
        pixel_data[483] = 3'b101; // x=3, y=12
        pixel_data[484] = 3'b101; // x=4, y=12
        pixel_data[485] = 3'b101; // x=5, y=12
        pixel_data[486] = 3'b101; // x=6, y=12
        pixel_data[487] = 3'b101; // x=7, y=12
        pixel_data[488] = 3'b101; // x=8, y=12
        pixel_data[489] = 3'b101; // x=9, y=12
        pixel_data[490] = 3'b101; // x=10, y=12
        pixel_data[491] = 3'b100; // x=11, y=12
        pixel_data[492] = 3'b100; // x=12, y=12
        pixel_data[493] = 3'b110; // x=13, y=12
        pixel_data[494] = 3'b110; // x=14, y=12
        pixel_data[495] = 3'b110; // x=15, y=12
        pixel_data[496] = 3'b110; // x=16, y=12
        pixel_data[497] = 3'b110; // x=17, y=12
        pixel_data[498] = 3'b110; // x=18, y=12
        pixel_data[499] = 3'b110; // x=19, y=12
        pixel_data[500] = 3'b110; // x=20, y=12
        pixel_data[501] = 3'b110; // x=21, y=12
        pixel_data[502] = 3'b110; // x=22, y=12
        pixel_data[503] = 3'b111; // x=23, y=12
        pixel_data[504] = 3'b110; // x=24, y=12
        pixel_data[505] = 3'b110; // x=25, y=12
        pixel_data[506] = 3'b111; // x=26, y=12
        pixel_data[507] = 3'b111; // x=27, y=12
        pixel_data[508] = 3'b110; // x=28, y=12
        pixel_data[509] = 3'b110; // x=29, y=12
        pixel_data[510] = 3'b101; // x=30, y=12
        pixel_data[511] = 3'b101; // x=31, y=12
        pixel_data[512] = 3'b101; // x=32, y=12
        pixel_data[513] = 3'b101; // x=33, y=12
        pixel_data[514] = 3'b101; // x=34, y=12
        pixel_data[515] = 3'b101; // x=35, y=12
        pixel_data[516] = 3'b101; // x=36, y=12
        pixel_data[517] = 3'b011; // x=37, y=12
        pixel_data[518] = 3'b001; // x=38, y=12
        pixel_data[519] = 3'b010; // x=39, y=12
        pixel_data[520] = 3'b010; // x=0, y=13
        pixel_data[521] = 3'b000; // x=1, y=13
        pixel_data[522] = 3'b100; // x=2, y=13
        pixel_data[523] = 3'b101; // x=3, y=13
        pixel_data[524] = 3'b101; // x=4, y=13
        pixel_data[525] = 3'b100; // x=5, y=13
        pixel_data[526] = 3'b101; // x=6, y=13
        pixel_data[527] = 3'b101; // x=7, y=13
        pixel_data[528] = 3'b101; // x=8, y=13
        pixel_data[529] = 3'b101; // x=9, y=13
        pixel_data[530] = 3'b101; // x=10, y=13
        pixel_data[531] = 3'b100; // x=11, y=13
        pixel_data[532] = 3'b101; // x=12, y=13
        pixel_data[533] = 3'b111; // x=13, y=13
        pixel_data[534] = 3'b110; // x=14, y=13
        pixel_data[535] = 3'b110; // x=15, y=13
        pixel_data[536] = 3'b110; // x=16, y=13
        pixel_data[537] = 3'b110; // x=17, y=13
        pixel_data[538] = 3'b110; // x=18, y=13
        pixel_data[539] = 3'b111; // x=19, y=13
        pixel_data[540] = 3'b111; // x=20, y=13
        pixel_data[541] = 3'b111; // x=21, y=13
        pixel_data[542] = 3'b111; // x=22, y=13
        pixel_data[543] = 3'b111; // x=23, y=13
        pixel_data[544] = 3'b111; // x=24, y=13
        pixel_data[545] = 3'b111; // x=25, y=13
        pixel_data[546] = 3'b111; // x=26, y=13
        pixel_data[547] = 3'b111; // x=27, y=13
        pixel_data[548] = 3'b111; // x=28, y=13
        pixel_data[549] = 3'b111; // x=29, y=13
        pixel_data[550] = 3'b111; // x=30, y=13
        pixel_data[551] = 3'b110; // x=31, y=13
        pixel_data[552] = 3'b110; // x=32, y=13
        pixel_data[553] = 3'b110; // x=33, y=13
        pixel_data[554] = 3'b101; // x=34, y=13
        pixel_data[555] = 3'b101; // x=35, y=13
        pixel_data[556] = 3'b101; // x=36, y=13
        pixel_data[557] = 3'b101; // x=37, y=13
        pixel_data[558] = 3'b000; // x=38, y=13
        pixel_data[559] = 3'b010; // x=39, y=13
        pixel_data[560] = 3'b001; // x=0, y=14
        pixel_data[561] = 3'b011; // x=1, y=14
        pixel_data[562] = 3'b101; // x=2, y=14
        pixel_data[563] = 3'b101; // x=3, y=14
        pixel_data[564] = 3'b101; // x=4, y=14
        pixel_data[565] = 3'b101; // x=5, y=14
        pixel_data[566] = 3'b101; // x=6, y=14
        pixel_data[567] = 3'b101; // x=7, y=14
        pixel_data[568] = 3'b101; // x=8, y=14
        pixel_data[569] = 3'b101; // x=9, y=14
        pixel_data[570] = 3'b101; // x=10, y=14
        pixel_data[571] = 3'b101; // x=11, y=14
        pixel_data[572] = 3'b111; // x=12, y=14
        pixel_data[573] = 3'b111; // x=13, y=14
        pixel_data[574] = 3'b110; // x=14, y=14
        pixel_data[575] = 3'b110; // x=15, y=14
        pixel_data[576] = 3'b110; // x=16, y=14
        pixel_data[577] = 3'b110; // x=17, y=14
        pixel_data[578] = 3'b110; // x=18, y=14
        pixel_data[579] = 3'b111; // x=19, y=14
        pixel_data[580] = 3'b111; // x=20, y=14
        pixel_data[581] = 3'b111; // x=21, y=14
        pixel_data[582] = 3'b111; // x=22, y=14
        pixel_data[583] = 3'b111; // x=23, y=14
        pixel_data[584] = 3'b111; // x=24, y=14
        pixel_data[585] = 3'b111; // x=25, y=14
        pixel_data[586] = 3'b111; // x=26, y=14
        pixel_data[587] = 3'b111; // x=27, y=14
        pixel_data[588] = 3'b111; // x=28, y=14
        pixel_data[589] = 3'b111; // x=29, y=14
        pixel_data[590] = 3'b111; // x=30, y=14
        pixel_data[591] = 3'b111; // x=31, y=14
        pixel_data[592] = 3'b111; // x=32, y=14
        pixel_data[593] = 3'b111; // x=33, y=14
        pixel_data[594] = 3'b111; // x=34, y=14
        pixel_data[595] = 3'b110; // x=35, y=14
        pixel_data[596] = 3'b101; // x=36, y=14
        pixel_data[597] = 3'b101; // x=37, y=14
        pixel_data[598] = 3'b011; // x=38, y=14
        pixel_data[599] = 3'b011; // x=39, y=14
        pixel_data[600] = 3'b000; // x=0, y=15
        pixel_data[601] = 3'b100; // x=1, y=15
        pixel_data[602] = 3'b101; // x=2, y=15
        pixel_data[603] = 3'b101; // x=3, y=15
        pixel_data[604] = 3'b100; // x=4, y=15
        pixel_data[605] = 3'b101; // x=5, y=15
        pixel_data[606] = 3'b101; // x=6, y=15
        pixel_data[607] = 3'b100; // x=7, y=15
        pixel_data[608] = 3'b100; // x=8, y=15
        pixel_data[609] = 3'b100; // x=9, y=15
        pixel_data[610] = 3'b100; // x=10, y=15
        pixel_data[611] = 3'b101; // x=11, y=15
        pixel_data[612] = 3'b111; // x=12, y=15
        pixel_data[613] = 3'b110; // x=13, y=15
        pixel_data[614] = 3'b110; // x=14, y=15
        pixel_data[615] = 3'b110; // x=15, y=15
        pixel_data[616] = 3'b110; // x=16, y=15
        pixel_data[617] = 3'b110; // x=17, y=15
        pixel_data[618] = 3'b111; // x=18, y=15
        pixel_data[619] = 3'b111; // x=19, y=15
        pixel_data[620] = 3'b111; // x=20, y=15
        pixel_data[621] = 3'b111; // x=21, y=15
        pixel_data[622] = 3'b111; // x=22, y=15
        pixel_data[623] = 3'b110; // x=23, y=15
        pixel_data[624] = 3'b111; // x=24, y=15
        pixel_data[625] = 3'b111; // x=25, y=15
        pixel_data[626] = 3'b111; // x=26, y=15
        pixel_data[627] = 3'b111; // x=27, y=15
        pixel_data[628] = 3'b111; // x=28, y=15
        pixel_data[629] = 3'b111; // x=29, y=15
        pixel_data[630] = 3'b111; // x=30, y=15
        pixel_data[631] = 3'b111; // x=31, y=15
        pixel_data[632] = 3'b111; // x=32, y=15
        pixel_data[633] = 3'b111; // x=33, y=15
        pixel_data[634] = 3'b111; // x=34, y=15
        pixel_data[635] = 3'b110; // x=35, y=15
        pixel_data[636] = 3'b100; // x=36, y=15
        pixel_data[637] = 3'b101; // x=37, y=15
        pixel_data[638] = 3'b100; // x=38, y=15
        pixel_data[639] = 3'b001; // x=39, y=15
        pixel_data[640] = 3'b000; // x=0, y=16
        pixel_data[641] = 3'b100; // x=1, y=16
        pixel_data[642] = 3'b101; // x=2, y=16
        pixel_data[643] = 3'b101; // x=3, y=16
        pixel_data[644] = 3'b101; // x=4, y=16
        pixel_data[645] = 3'b101; // x=5, y=16
        pixel_data[646] = 3'b100; // x=6, y=16
        pixel_data[647] = 3'b100; // x=7, y=16
        pixel_data[648] = 3'b100; // x=8, y=16
        pixel_data[649] = 3'b100; // x=9, y=16
        pixel_data[650] = 3'b100; // x=10, y=16
        pixel_data[651] = 3'b110; // x=11, y=16
        pixel_data[652] = 3'b111; // x=12, y=16
        pixel_data[653] = 3'b110; // x=13, y=16
        pixel_data[654] = 3'b110; // x=14, y=16
        pixel_data[655] = 3'b110; // x=15, y=16
        pixel_data[656] = 3'b110; // x=16, y=16
        pixel_data[657] = 3'b110; // x=17, y=16
        pixel_data[658] = 3'b111; // x=18, y=16
        pixel_data[659] = 3'b111; // x=19, y=16
        pixel_data[660] = 3'b111; // x=20, y=16
        pixel_data[661] = 3'b111; // x=21, y=16
        pixel_data[662] = 3'b111; // x=22, y=16
        pixel_data[663] = 3'b110; // x=23, y=16
        pixel_data[664] = 3'b111; // x=24, y=16
        pixel_data[665] = 3'b111; // x=25, y=16
        pixel_data[666] = 3'b111; // x=26, y=16
        pixel_data[667] = 3'b111; // x=27, y=16
        pixel_data[668] = 3'b111; // x=28, y=16
        pixel_data[669] = 3'b111; // x=29, y=16
        pixel_data[670] = 3'b111; // x=30, y=16
        pixel_data[671] = 3'b111; // x=31, y=16
        pixel_data[672] = 3'b111; // x=32, y=16
        pixel_data[673] = 3'b111; // x=33, y=16
        pixel_data[674] = 3'b111; // x=34, y=16
        pixel_data[675] = 3'b110; // x=35, y=16
        pixel_data[676] = 3'b100; // x=36, y=16
        pixel_data[677] = 3'b101; // x=37, y=16
        pixel_data[678] = 3'b100; // x=38, y=16
        pixel_data[679] = 3'b000; // x=39, y=16
        pixel_data[680] = 3'b000; // x=0, y=17
        pixel_data[681] = 3'b100; // x=1, y=17
        pixel_data[682] = 3'b101; // x=2, y=17
        pixel_data[683] = 3'b101; // x=3, y=17
        pixel_data[684] = 3'b101; // x=4, y=17
        pixel_data[685] = 3'b100; // x=5, y=17
        pixel_data[686] = 3'b100; // x=6, y=17
        pixel_data[687] = 3'b100; // x=7, y=17
        pixel_data[688] = 3'b100; // x=8, y=17
        pixel_data[689] = 3'b100; // x=9, y=17
        pixel_data[690] = 3'b100; // x=10, y=17
        pixel_data[691] = 3'b110; // x=11, y=17
        pixel_data[692] = 3'b111; // x=12, y=17
        pixel_data[693] = 3'b110; // x=13, y=17
        pixel_data[694] = 3'b110; // x=14, y=17
        pixel_data[695] = 3'b110; // x=15, y=17
        pixel_data[696] = 3'b110; // x=16, y=17
        pixel_data[697] = 3'b110; // x=17, y=17
        pixel_data[698] = 3'b111; // x=18, y=17
        pixel_data[699] = 3'b111; // x=19, y=17
        pixel_data[700] = 3'b111; // x=20, y=17
        pixel_data[701] = 3'b111; // x=21, y=17
        pixel_data[702] = 3'b111; // x=22, y=17
        pixel_data[703] = 3'b110; // x=23, y=17
        pixel_data[704] = 3'b111; // x=24, y=17
        pixel_data[705] = 3'b111; // x=25, y=17
        pixel_data[706] = 3'b111; // x=26, y=17
        pixel_data[707] = 3'b111; // x=27, y=17
        pixel_data[708] = 3'b111; // x=28, y=17
        pixel_data[709] = 3'b111; // x=29, y=17
        pixel_data[710] = 3'b111; // x=30, y=17
        pixel_data[711] = 3'b111; // x=31, y=17
        pixel_data[712] = 3'b111; // x=32, y=17
        pixel_data[713] = 3'b111; // x=33, y=17
        pixel_data[714] = 3'b111; // x=34, y=17
        pixel_data[715] = 3'b110; // x=35, y=17
        pixel_data[716] = 3'b100; // x=36, y=17
        pixel_data[717] = 3'b101; // x=37, y=17
        pixel_data[718] = 3'b101; // x=38, y=17
        pixel_data[719] = 3'b000; // x=39, y=17
        pixel_data[720] = 3'b000; // x=0, y=18
        pixel_data[721] = 3'b101; // x=1, y=18
        pixel_data[722] = 3'b101; // x=2, y=18
        pixel_data[723] = 3'b101; // x=3, y=18
        pixel_data[724] = 3'b100; // x=4, y=18
        pixel_data[725] = 3'b100; // x=5, y=18
        pixel_data[726] = 3'b100; // x=6, y=18
        pixel_data[727] = 3'b100; // x=7, y=18
        pixel_data[728] = 3'b100; // x=8, y=18
        pixel_data[729] = 3'b100; // x=9, y=18
        pixel_data[730] = 3'b101; // x=10, y=18
        pixel_data[731] = 3'b111; // x=11, y=18
        pixel_data[732] = 3'b111; // x=12, y=18
        pixel_data[733] = 3'b110; // x=13, y=18
        pixel_data[734] = 3'b110; // x=14, y=18
        pixel_data[735] = 3'b110; // x=15, y=18
        pixel_data[736] = 3'b110; // x=16, y=18
        pixel_data[737] = 3'b110; // x=17, y=18
        pixel_data[738] = 3'b111; // x=18, y=18
        pixel_data[739] = 3'b111; // x=19, y=18
        pixel_data[740] = 3'b111; // x=20, y=18
        pixel_data[741] = 3'b111; // x=21, y=18
        pixel_data[742] = 3'b111; // x=22, y=18
        pixel_data[743] = 3'b110; // x=23, y=18
        pixel_data[744] = 3'b111; // x=24, y=18
        pixel_data[745] = 3'b111; // x=25, y=18
        pixel_data[746] = 3'b111; // x=26, y=18
        pixel_data[747] = 3'b111; // x=27, y=18
        pixel_data[748] = 3'b111; // x=28, y=18
        pixel_data[749] = 3'b111; // x=29, y=18
        pixel_data[750] = 3'b111; // x=30, y=18
        pixel_data[751] = 3'b111; // x=31, y=18
        pixel_data[752] = 3'b111; // x=32, y=18
        pixel_data[753] = 3'b111; // x=33, y=18
        pixel_data[754] = 3'b111; // x=34, y=18
        pixel_data[755] = 3'b110; // x=35, y=18
        pixel_data[756] = 3'b100; // x=36, y=18
        pixel_data[757] = 3'b101; // x=37, y=18
        pixel_data[758] = 3'b101; // x=38, y=18
        pixel_data[759] = 3'b001; // x=39, y=18
        pixel_data[760] = 3'b000; // x=0, y=19
        pixel_data[761] = 3'b101; // x=1, y=19
        pixel_data[762] = 3'b101; // x=2, y=19
        pixel_data[763] = 3'b101; // x=3, y=19
        pixel_data[764] = 3'b100; // x=4, y=19
        pixel_data[765] = 3'b100; // x=5, y=19
        pixel_data[766] = 3'b100; // x=6, y=19
        pixel_data[767] = 3'b100; // x=7, y=19
        pixel_data[768] = 3'b100; // x=8, y=19
        pixel_data[769] = 3'b100; // x=9, y=19
        pixel_data[770] = 3'b101; // x=10, y=19
        pixel_data[771] = 3'b111; // x=11, y=19
        pixel_data[772] = 3'b111; // x=12, y=19
        pixel_data[773] = 3'b110; // x=13, y=19
        pixel_data[774] = 3'b110; // x=14, y=19
        pixel_data[775] = 3'b110; // x=15, y=19
        pixel_data[776] = 3'b110; // x=16, y=19
        pixel_data[777] = 3'b110; // x=17, y=19
        pixel_data[778] = 3'b111; // x=18, y=19
        pixel_data[779] = 3'b111; // x=19, y=19
        pixel_data[780] = 3'b111; // x=20, y=19
        pixel_data[781] = 3'b111; // x=21, y=19
        pixel_data[782] = 3'b111; // x=22, y=19
        pixel_data[783] = 3'b110; // x=23, y=19
        pixel_data[784] = 3'b111; // x=24, y=19
        pixel_data[785] = 3'b111; // x=25, y=19
        pixel_data[786] = 3'b111; // x=26, y=19
        pixel_data[787] = 3'b111; // x=27, y=19
        pixel_data[788] = 3'b111; // x=28, y=19
        pixel_data[789] = 3'b111; // x=29, y=19
        pixel_data[790] = 3'b111; // x=30, y=19
        pixel_data[791] = 3'b111; // x=31, y=19
        pixel_data[792] = 3'b111; // x=32, y=19
        pixel_data[793] = 3'b111; // x=33, y=19
        pixel_data[794] = 3'b111; // x=34, y=19
        pixel_data[795] = 3'b110; // x=35, y=19
        pixel_data[796] = 3'b100; // x=36, y=19
        pixel_data[797] = 3'b101; // x=37, y=19
        pixel_data[798] = 3'b101; // x=38, y=19
        pixel_data[799] = 3'b011; // x=39, y=19
        pixel_data[800] = 3'b000; // x=0, y=20
        pixel_data[801] = 3'b101; // x=1, y=20
        pixel_data[802] = 3'b101; // x=2, y=20
        pixel_data[803] = 3'b101; // x=3, y=20
        pixel_data[804] = 3'b100; // x=4, y=20
        pixel_data[805] = 3'b100; // x=5, y=20
        pixel_data[806] = 3'b100; // x=6, y=20
        pixel_data[807] = 3'b100; // x=7, y=20
        pixel_data[808] = 3'b100; // x=8, y=20
        pixel_data[809] = 3'b100; // x=9, y=20
        pixel_data[810] = 3'b101; // x=10, y=20
        pixel_data[811] = 3'b111; // x=11, y=20
        pixel_data[812] = 3'b111; // x=12, y=20
        pixel_data[813] = 3'b110; // x=13, y=20
        pixel_data[814] = 3'b110; // x=14, y=20
        pixel_data[815] = 3'b110; // x=15, y=20
        pixel_data[816] = 3'b110; // x=16, y=20
        pixel_data[817] = 3'b110; // x=17, y=20
        pixel_data[818] = 3'b111; // x=18, y=20
        pixel_data[819] = 3'b111; // x=19, y=20
        pixel_data[820] = 3'b111; // x=20, y=20
        pixel_data[821] = 3'b111; // x=21, y=20
        pixel_data[822] = 3'b111; // x=22, y=20
        pixel_data[823] = 3'b110; // x=23, y=20
        pixel_data[824] = 3'b111; // x=24, y=20
        pixel_data[825] = 3'b111; // x=25, y=20
        pixel_data[826] = 3'b111; // x=26, y=20
        pixel_data[827] = 3'b111; // x=27, y=20
        pixel_data[828] = 3'b111; // x=28, y=20
        pixel_data[829] = 3'b111; // x=29, y=20
        pixel_data[830] = 3'b111; // x=30, y=20
        pixel_data[831] = 3'b111; // x=31, y=20
        pixel_data[832] = 3'b111; // x=32, y=20
        pixel_data[833] = 3'b111; // x=33, y=20
        pixel_data[834] = 3'b111; // x=34, y=20
        pixel_data[835] = 3'b110; // x=35, y=20
        pixel_data[836] = 3'b100; // x=36, y=20
        pixel_data[837] = 3'b101; // x=37, y=20
        pixel_data[838] = 3'b101; // x=38, y=20
        pixel_data[839] = 3'b010; // x=39, y=20
        pixel_data[840] = 3'b000; // x=0, y=21
        pixel_data[841] = 3'b100; // x=1, y=21
        pixel_data[842] = 3'b101; // x=2, y=21
        pixel_data[843] = 3'b101; // x=3, y=21
        pixel_data[844] = 3'b100; // x=4, y=21
        pixel_data[845] = 3'b100; // x=5, y=21
        pixel_data[846] = 3'b100; // x=6, y=21
        pixel_data[847] = 3'b100; // x=7, y=21
        pixel_data[848] = 3'b100; // x=8, y=21
        pixel_data[849] = 3'b100; // x=9, y=21
        pixel_data[850] = 3'b100; // x=10, y=21
        pixel_data[851] = 3'b110; // x=11, y=21
        pixel_data[852] = 3'b111; // x=12, y=21
        pixel_data[853] = 3'b110; // x=13, y=21
        pixel_data[854] = 3'b110; // x=14, y=21
        pixel_data[855] = 3'b110; // x=15, y=21
        pixel_data[856] = 3'b110; // x=16, y=21
        pixel_data[857] = 3'b110; // x=17, y=21
        pixel_data[858] = 3'b111; // x=18, y=21
        pixel_data[859] = 3'b111; // x=19, y=21
        pixel_data[860] = 3'b111; // x=20, y=21
        pixel_data[861] = 3'b111; // x=21, y=21
        pixel_data[862] = 3'b111; // x=22, y=21
        pixel_data[863] = 3'b110; // x=23, y=21
        pixel_data[864] = 3'b111; // x=24, y=21
        pixel_data[865] = 3'b111; // x=25, y=21
        pixel_data[866] = 3'b111; // x=26, y=21
        pixel_data[867] = 3'b111; // x=27, y=21
        pixel_data[868] = 3'b111; // x=28, y=21
        pixel_data[869] = 3'b111; // x=29, y=21
        pixel_data[870] = 3'b111; // x=30, y=21
        pixel_data[871] = 3'b111; // x=31, y=21
        pixel_data[872] = 3'b111; // x=32, y=21
        pixel_data[873] = 3'b111; // x=33, y=21
        pixel_data[874] = 3'b111; // x=34, y=21
        pixel_data[875] = 3'b110; // x=35, y=21
        pixel_data[876] = 3'b100; // x=36, y=21
        pixel_data[877] = 3'b101; // x=37, y=21
        pixel_data[878] = 3'b101; // x=38, y=21
        pixel_data[879] = 3'b000; // x=39, y=21
        pixel_data[880] = 3'b000; // x=0, y=22
        pixel_data[881] = 3'b100; // x=1, y=22
        pixel_data[882] = 3'b101; // x=2, y=22
        pixel_data[883] = 3'b101; // x=3, y=22
        pixel_data[884] = 3'b100; // x=4, y=22
        pixel_data[885] = 3'b100; // x=5, y=22
        pixel_data[886] = 3'b100; // x=6, y=22
        pixel_data[887] = 3'b100; // x=7, y=22
        pixel_data[888] = 3'b100; // x=8, y=22
        pixel_data[889] = 3'b100; // x=9, y=22
        pixel_data[890] = 3'b100; // x=10, y=22
        pixel_data[891] = 3'b110; // x=11, y=22
        pixel_data[892] = 3'b111; // x=12, y=22
        pixel_data[893] = 3'b110; // x=13, y=22
        pixel_data[894] = 3'b110; // x=14, y=22
        pixel_data[895] = 3'b110; // x=15, y=22
        pixel_data[896] = 3'b110; // x=16, y=22
        pixel_data[897] = 3'b110; // x=17, y=22
        pixel_data[898] = 3'b111; // x=18, y=22
        pixel_data[899] = 3'b111; // x=19, y=22
        pixel_data[900] = 3'b111; // x=20, y=22
        pixel_data[901] = 3'b111; // x=21, y=22
        pixel_data[902] = 3'b111; // x=22, y=22
        pixel_data[903] = 3'b110; // x=23, y=22
        pixel_data[904] = 3'b111; // x=24, y=22
        pixel_data[905] = 3'b111; // x=25, y=22
        pixel_data[906] = 3'b111; // x=26, y=22
        pixel_data[907] = 3'b111; // x=27, y=22
        pixel_data[908] = 3'b111; // x=28, y=22
        pixel_data[909] = 3'b111; // x=29, y=22
        pixel_data[910] = 3'b111; // x=30, y=22
        pixel_data[911] = 3'b111; // x=31, y=22
        pixel_data[912] = 3'b111; // x=32, y=22
        pixel_data[913] = 3'b111; // x=33, y=22
        pixel_data[914] = 3'b111; // x=34, y=22
        pixel_data[915] = 3'b110; // x=35, y=22
        pixel_data[916] = 3'b100; // x=36, y=22
        pixel_data[917] = 3'b101; // x=37, y=22
        pixel_data[918] = 3'b100; // x=38, y=22
        pixel_data[919] = 3'b000; // x=39, y=22
        pixel_data[920] = 3'b000; // x=0, y=23
        pixel_data[921] = 3'b100; // x=1, y=23
        pixel_data[922] = 3'b101; // x=2, y=23
        pixel_data[923] = 3'b101; // x=3, y=23
        pixel_data[924] = 3'b101; // x=4, y=23
        pixel_data[925] = 3'b101; // x=5, y=23
        pixel_data[926] = 3'b101; // x=6, y=23
        pixel_data[927] = 3'b101; // x=7, y=23
        pixel_data[928] = 3'b101; // x=8, y=23
        pixel_data[929] = 3'b101; // x=9, y=23
        pixel_data[930] = 3'b100; // x=10, y=23
        pixel_data[931] = 3'b101; // x=11, y=23
        pixel_data[932] = 3'b111; // x=12, y=23
        pixel_data[933] = 3'b110; // x=13, y=23
        pixel_data[934] = 3'b110; // x=14, y=23
        pixel_data[935] = 3'b110; // x=15, y=23
        pixel_data[936] = 3'b110; // x=16, y=23
        pixel_data[937] = 3'b110; // x=17, y=23
        pixel_data[938] = 3'b111; // x=18, y=23
        pixel_data[939] = 3'b111; // x=19, y=23
        pixel_data[940] = 3'b110; // x=20, y=23
        pixel_data[941] = 3'b111; // x=21, y=23
        pixel_data[942] = 3'b111; // x=22, y=23
        pixel_data[943] = 3'b110; // x=23, y=23
        pixel_data[944] = 3'b111; // x=24, y=23
        pixel_data[945] = 3'b111; // x=25, y=23
        pixel_data[946] = 3'b111; // x=26, y=23
        pixel_data[947] = 3'b111; // x=27, y=23
        pixel_data[948] = 3'b111; // x=28, y=23
        pixel_data[949] = 3'b111; // x=29, y=23
        pixel_data[950] = 3'b111; // x=30, y=23
        pixel_data[951] = 3'b111; // x=31, y=23
        pixel_data[952] = 3'b111; // x=32, y=23
        pixel_data[953] = 3'b111; // x=33, y=23
        pixel_data[954] = 3'b111; // x=34, y=23
        pixel_data[955] = 3'b110; // x=35, y=23
        pixel_data[956] = 3'b100; // x=36, y=23
        pixel_data[957] = 3'b101; // x=37, y=23
        pixel_data[958] = 3'b100; // x=38, y=23
        pixel_data[959] = 3'b000; // x=39, y=23
        pixel_data[960] = 3'b010; // x=0, y=24
        pixel_data[961] = 3'b011; // x=1, y=24
        pixel_data[962] = 3'b101; // x=2, y=24
        pixel_data[963] = 3'b101; // x=3, y=24
        pixel_data[964] = 3'b101; // x=4, y=24
        pixel_data[965] = 3'b101; // x=5, y=24
        pixel_data[966] = 3'b101; // x=6, y=24
        pixel_data[967] = 3'b101; // x=7, y=24
        pixel_data[968] = 3'b101; // x=8, y=24
        pixel_data[969] = 3'b101; // x=9, y=24
        pixel_data[970] = 3'b101; // x=10, y=24
        pixel_data[971] = 3'b101; // x=11, y=24
        pixel_data[972] = 3'b110; // x=12, y=24
        pixel_data[973] = 3'b111; // x=13, y=24
        pixel_data[974] = 3'b110; // x=14, y=24
        pixel_data[975] = 3'b110; // x=15, y=24
        pixel_data[976] = 3'b110; // x=16, y=24
        pixel_data[977] = 3'b110; // x=17, y=24
        pixel_data[978] = 3'b110; // x=18, y=24
        pixel_data[979] = 3'b111; // x=19, y=24
        pixel_data[980] = 3'b111; // x=20, y=24
        pixel_data[981] = 3'b111; // x=21, y=24
        pixel_data[982] = 3'b111; // x=22, y=24
        pixel_data[983] = 3'b111; // x=23, y=24
        pixel_data[984] = 3'b111; // x=24, y=24
        pixel_data[985] = 3'b111; // x=25, y=24
        pixel_data[986] = 3'b111; // x=26, y=24
        pixel_data[987] = 3'b111; // x=27, y=24
        pixel_data[988] = 3'b111; // x=28, y=24
        pixel_data[989] = 3'b111; // x=29, y=24
        pixel_data[990] = 3'b111; // x=30, y=24
        pixel_data[991] = 3'b111; // x=31, y=24
        pixel_data[992] = 3'b111; // x=32, y=24
        pixel_data[993] = 3'b111; // x=33, y=24
        pixel_data[994] = 3'b111; // x=34, y=24
        pixel_data[995] = 3'b110; // x=35, y=24
        pixel_data[996] = 3'b101; // x=36, y=24
        pixel_data[997] = 3'b101; // x=37, y=24
        pixel_data[998] = 3'b011; // x=38, y=24
        pixel_data[999] = 3'b001; // x=39, y=24
        pixel_data[1000] = 3'b010; // x=0, y=25
        pixel_data[1001] = 3'b000; // x=1, y=25
        pixel_data[1002] = 3'b100; // x=2, y=25
        pixel_data[1003] = 3'b101; // x=3, y=25
        pixel_data[1004] = 3'b101; // x=4, y=25
        pixel_data[1005] = 3'b100; // x=5, y=25
        pixel_data[1006] = 3'b100; // x=6, y=25
        pixel_data[1007] = 3'b100; // x=7, y=25
        pixel_data[1008] = 3'b100; // x=8, y=25
        pixel_data[1009] = 3'b100; // x=9, y=25
        pixel_data[1010] = 3'b100; // x=10, y=25
        pixel_data[1011] = 3'b100; // x=11, y=25
        pixel_data[1012] = 3'b101; // x=12, y=25
        pixel_data[1013] = 3'b111; // x=13, y=25
        pixel_data[1014] = 3'b110; // x=14, y=25
        pixel_data[1015] = 3'b110; // x=15, y=25
        pixel_data[1016] = 3'b110; // x=16, y=25
        pixel_data[1017] = 3'b110; // x=17, y=25
        pixel_data[1018] = 3'b110; // x=18, y=25
        pixel_data[1019] = 3'b111; // x=19, y=25
        pixel_data[1020] = 3'b111; // x=20, y=25
        pixel_data[1021] = 3'b111; // x=21, y=25
        pixel_data[1022] = 3'b111; // x=22, y=25
        pixel_data[1023] = 3'b111; // x=23, y=25
        pixel_data[1024] = 3'b111; // x=24, y=25
        pixel_data[1025] = 3'b111; // x=25, y=25
        pixel_data[1026] = 3'b111; // x=26, y=25
        pixel_data[1027] = 3'b111; // x=27, y=25
        pixel_data[1028] = 3'b111; // x=28, y=25
        pixel_data[1029] = 3'b111; // x=29, y=25
        pixel_data[1030] = 3'b111; // x=30, y=25
        pixel_data[1031] = 3'b110; // x=31, y=25
        pixel_data[1032] = 3'b110; // x=32, y=25
        pixel_data[1033] = 3'b101; // x=33, y=25
        pixel_data[1034] = 3'b101; // x=34, y=25
        pixel_data[1035] = 3'b101; // x=35, y=25
        pixel_data[1036] = 3'b101; // x=36, y=25
        pixel_data[1037] = 3'b101; // x=37, y=25
        pixel_data[1038] = 3'b001; // x=38, y=25
        pixel_data[1039] = 3'b011; // x=39, y=25
        pixel_data[1040] = 3'b010; // x=0, y=26
        pixel_data[1041] = 3'b001; // x=1, y=26
        pixel_data[1042] = 3'b011; // x=2, y=26
        pixel_data[1043] = 3'b101; // x=3, y=26
        pixel_data[1044] = 3'b101; // x=4, y=26
        pixel_data[1045] = 3'b101; // x=5, y=26
        pixel_data[1046] = 3'b101; // x=6, y=26
        pixel_data[1047] = 3'b101; // x=7, y=26
        pixel_data[1048] = 3'b101; // x=8, y=26
        pixel_data[1049] = 3'b101; // x=9, y=26
        pixel_data[1050] = 3'b101; // x=10, y=26
        pixel_data[1051] = 3'b101; // x=11, y=26
        pixel_data[1052] = 3'b101; // x=12, y=26
        pixel_data[1053] = 3'b110; // x=13, y=26
        pixel_data[1054] = 3'b110; // x=14, y=26
        pixel_data[1055] = 3'b110; // x=15, y=26
        pixel_data[1056] = 3'b110; // x=16, y=26
        pixel_data[1057] = 3'b110; // x=17, y=26
        pixel_data[1058] = 3'b110; // x=18, y=26
        pixel_data[1059] = 3'b110; // x=19, y=26
        pixel_data[1060] = 3'b111; // x=20, y=26
        pixel_data[1061] = 3'b111; // x=21, y=26
        pixel_data[1062] = 3'b111; // x=22, y=26
        pixel_data[1063] = 3'b111; // x=23, y=26
        pixel_data[1064] = 3'b110; // x=24, y=26
        pixel_data[1065] = 3'b111; // x=25, y=26
        pixel_data[1066] = 3'b111; // x=26, y=26
        pixel_data[1067] = 3'b111; // x=27, y=26
        pixel_data[1068] = 3'b111; // x=28, y=26
        pixel_data[1069] = 3'b111; // x=29, y=26
        pixel_data[1070] = 3'b110; // x=30, y=26
        pixel_data[1071] = 3'b101; // x=31, y=26
        pixel_data[1072] = 3'b101; // x=32, y=26
        pixel_data[1073] = 3'b101; // x=33, y=26
        pixel_data[1074] = 3'b101; // x=34, y=26
        pixel_data[1075] = 3'b101; // x=35, y=26
        pixel_data[1076] = 3'b101; // x=36, y=26
        pixel_data[1077] = 3'b011; // x=37, y=26
        pixel_data[1078] = 3'b011; // x=38, y=26
        pixel_data[1079] = 3'b011; // x=39, y=26
        pixel_data[1080] = 3'b010; // x=0, y=27
        pixel_data[1081] = 3'b010; // x=1, y=27
        pixel_data[1082] = 3'b001; // x=2, y=27
        pixel_data[1083] = 3'b011; // x=3, y=27
        pixel_data[1084] = 3'b100; // x=4, y=27
        pixel_data[1085] = 3'b101; // x=5, y=27
        pixel_data[1086] = 3'b101; // x=6, y=27
        pixel_data[1087] = 3'b101; // x=7, y=27
        pixel_data[1088] = 3'b101; // x=8, y=27
        pixel_data[1089] = 3'b101; // x=9, y=27
        pixel_data[1090] = 3'b101; // x=10, y=27
        pixel_data[1091] = 3'b101; // x=11, y=27
        pixel_data[1092] = 3'b101; // x=12, y=27
        pixel_data[1093] = 3'b101; // x=13, y=27
        pixel_data[1094] = 3'b101; // x=14, y=27
        pixel_data[1095] = 3'b110; // x=15, y=27
        pixel_data[1096] = 3'b110; // x=16, y=27
        pixel_data[1097] = 3'b110; // x=17, y=27
        pixel_data[1098] = 3'b110; // x=18, y=27
        pixel_data[1099] = 3'b110; // x=19, y=27
        pixel_data[1100] = 3'b110; // x=20, y=27
        pixel_data[1101] = 3'b110; // x=21, y=27
        pixel_data[1102] = 3'b110; // x=22, y=27
        pixel_data[1103] = 3'b110; // x=23, y=27
        pixel_data[1104] = 3'b110; // x=24, y=27
        pixel_data[1105] = 3'b110; // x=25, y=27
        pixel_data[1106] = 3'b110; // x=26, y=27
        pixel_data[1107] = 3'b110; // x=27, y=27
        pixel_data[1108] = 3'b110; // x=28, y=27
        pixel_data[1109] = 3'b110; // x=29, y=27
        pixel_data[1110] = 3'b101; // x=30, y=27
        pixel_data[1111] = 3'b101; // x=31, y=27
        pixel_data[1112] = 3'b101; // x=32, y=27
        pixel_data[1113] = 3'b100; // x=33, y=27
        pixel_data[1114] = 3'b100; // x=34, y=27
        pixel_data[1115] = 3'b100; // x=35, y=27
        pixel_data[1116] = 3'b011; // x=36, y=27
        pixel_data[1117] = 3'b011; // x=37, y=27
        pixel_data[1118] = 3'b011; // x=38, y=27
        pixel_data[1119] = 3'b010; // x=39, y=27
        pixel_data[1120] = 3'b010; // x=0, y=28
        pixel_data[1121] = 3'b010; // x=1, y=28
        pixel_data[1122] = 3'b010; // x=2, y=28
        pixel_data[1123] = 3'b011; // x=3, y=28
        pixel_data[1124] = 3'b010; // x=4, y=28
        pixel_data[1125] = 3'b000; // x=5, y=28
        pixel_data[1126] = 3'b001; // x=6, y=28
        pixel_data[1127] = 3'b010; // x=7, y=28
        pixel_data[1128] = 3'b011; // x=8, y=28
        pixel_data[1129] = 3'b011; // x=9, y=28
        pixel_data[1130] = 3'b011; // x=10, y=28
        pixel_data[1131] = 3'b011; // x=11, y=28
        pixel_data[1132] = 3'b011; // x=12, y=28
        pixel_data[1133] = 3'b011; // x=13, y=28
        pixel_data[1134] = 3'b011; // x=14, y=28
        pixel_data[1135] = 3'b101; // x=15, y=28
        pixel_data[1136] = 3'b101; // x=16, y=28
        pixel_data[1137] = 3'b000; // x=17, y=28
        pixel_data[1138] = 3'b000; // x=18, y=28
        pixel_data[1139] = 3'b000; // x=19, y=28
        pixel_data[1140] = 3'b000; // x=20, y=28
        pixel_data[1141] = 3'b000; // x=21, y=28
        pixel_data[1142] = 3'b011; // x=22, y=28
        pixel_data[1143] = 3'b100; // x=23, y=28
        pixel_data[1144] = 3'b000; // x=24, y=28
        pixel_data[1145] = 3'b011; // x=25, y=28
        pixel_data[1146] = 3'b100; // x=26, y=28
        pixel_data[1147] = 3'b000; // x=27, y=28
        pixel_data[1148] = 3'b000; // x=28, y=28
        pixel_data[1149] = 3'b000; // x=29, y=28
        pixel_data[1150] = 3'b000; // x=30, y=28
        pixel_data[1151] = 3'b000; // x=31, y=28
        pixel_data[1152] = 3'b000; // x=32, y=28
        pixel_data[1153] = 3'b000; // x=33, y=28
        pixel_data[1154] = 3'b000; // x=34, y=28
        pixel_data[1155] = 3'b000; // x=35, y=28
        pixel_data[1156] = 3'b011; // x=36, y=28
        pixel_data[1157] = 3'b011; // x=37, y=28
        pixel_data[1158] = 3'b010; // x=38, y=28
        pixel_data[1159] = 3'b010; // x=39, y=28
        pixel_data[1160] = 3'b010; // x=0, y=29
        pixel_data[1161] = 3'b010; // x=1, y=29
        pixel_data[1162] = 3'b011; // x=2, y=29
        pixel_data[1163] = 3'b010; // x=3, y=29
        pixel_data[1164] = 3'b010; // x=4, y=29
        pixel_data[1165] = 3'b010; // x=5, y=29
        pixel_data[1166] = 3'b010; // x=6, y=29
        pixel_data[1167] = 3'b010; // x=7, y=29
        pixel_data[1168] = 3'b010; // x=8, y=29
        pixel_data[1169] = 3'b010; // x=9, y=29
        pixel_data[1170] = 3'b010; // x=10, y=29
        pixel_data[1171] = 3'b010; // x=11, y=29
        pixel_data[1172] = 3'b010; // x=12, y=29
        pixel_data[1173] = 3'b010; // x=13, y=29
        pixel_data[1174] = 3'b001; // x=14, y=29
        pixel_data[1175] = 3'b100; // x=15, y=29
        pixel_data[1176] = 3'b100; // x=16, y=29
        pixel_data[1177] = 3'b000; // x=17, y=29
        pixel_data[1178] = 3'b010; // x=18, y=29
        pixel_data[1179] = 3'b010; // x=19, y=29
        pixel_data[1180] = 3'b001; // x=20, y=29
        pixel_data[1181] = 3'b001; // x=21, y=29
        pixel_data[1182] = 3'b000; // x=22, y=29
        pixel_data[1183] = 3'b000; // x=23, y=29
        pixel_data[1184] = 3'b010; // x=24, y=29
        pixel_data[1185] = 3'b001; // x=25, y=29
        pixel_data[1186] = 3'b000; // x=26, y=29
        pixel_data[1187] = 3'b001; // x=27, y=29
        pixel_data[1188] = 3'b010; // x=28, y=29
        pixel_data[1189] = 3'b010; // x=29, y=29
        pixel_data[1190] = 3'b010; // x=30, y=29
        pixel_data[1191] = 3'b010; // x=31, y=29
        pixel_data[1192] = 3'b010; // x=32, y=29
        pixel_data[1193] = 3'b010; // x=33, y=29
        pixel_data[1194] = 3'b010; // x=34, y=29
        pixel_data[1195] = 3'b011; // x=35, y=29
        pixel_data[1196] = 3'b010; // x=36, y=29
        pixel_data[1197] = 3'b010; // x=37, y=29
        pixel_data[1198] = 3'b010; // x=38, y=29
        pixel_data[1199] = 3'b010; // x=39, y=29
        pixel_data[1200] = 3'b010; // x=0, y=30
        pixel_data[1201] = 3'b010; // x=1, y=30
        pixel_data[1202] = 3'b010; // x=2, y=30
        pixel_data[1203] = 3'b010; // x=3, y=30
        pixel_data[1204] = 3'b010; // x=4, y=30
        pixel_data[1205] = 3'b010; // x=5, y=30
        pixel_data[1206] = 3'b010; // x=6, y=30
        pixel_data[1207] = 3'b010; // x=7, y=30
        pixel_data[1208] = 3'b011; // x=8, y=30
        pixel_data[1209] = 3'b010; // x=9, y=30
        pixel_data[1210] = 3'b010; // x=10, y=30
        pixel_data[1211] = 3'b010; // x=11, y=30
        pixel_data[1212] = 3'b011; // x=12, y=30
        pixel_data[1213] = 3'b011; // x=13, y=30
        pixel_data[1214] = 3'b010; // x=14, y=30
        pixel_data[1215] = 3'b001; // x=15, y=30
        pixel_data[1216] = 3'b000; // x=16, y=30
        pixel_data[1217] = 3'b010; // x=17, y=30
        pixel_data[1218] = 3'b010; // x=18, y=30
        pixel_data[1219] = 3'b011; // x=19, y=30
        pixel_data[1220] = 3'b010; // x=20, y=30
        pixel_data[1221] = 3'b010; // x=21, y=30
        pixel_data[1222] = 3'b010; // x=22, y=30
        pixel_data[1223] = 3'b010; // x=23, y=30
        pixel_data[1224] = 3'b010; // x=24, y=30
        pixel_data[1225] = 3'b010; // x=25, y=30
        pixel_data[1226] = 3'b010; // x=26, y=30
        pixel_data[1227] = 3'b010; // x=27, y=30
        pixel_data[1228] = 3'b010; // x=28, y=30
        pixel_data[1229] = 3'b010; // x=29, y=30
        pixel_data[1230] = 3'b011; // x=30, y=30
        pixel_data[1231] = 3'b010; // x=31, y=30
        pixel_data[1232] = 3'b010; // x=32, y=30
        pixel_data[1233] = 3'b010; // x=33, y=30
        pixel_data[1234] = 3'b011; // x=34, y=30
        pixel_data[1235] = 3'b010; // x=35, y=30
        pixel_data[1236] = 3'b010; // x=36, y=30
        pixel_data[1237] = 3'b010; // x=37, y=30
        pixel_data[1238] = 3'b010; // x=38, y=30
        pixel_data[1239] = 3'b010; // x=39, y=30
        pixel_data[1240] = 3'b010; // x=0, y=31
        pixel_data[1241] = 3'b010; // x=1, y=31
        pixel_data[1242] = 3'b010; // x=2, y=31
        pixel_data[1243] = 3'b010; // x=3, y=31
        pixel_data[1244] = 3'b010; // x=4, y=31
        pixel_data[1245] = 3'b010; // x=5, y=31
        pixel_data[1246] = 3'b010; // x=6, y=31
        pixel_data[1247] = 3'b010; // x=7, y=31
        pixel_data[1248] = 3'b010; // x=8, y=31
        pixel_data[1249] = 3'b011; // x=9, y=31
        pixel_data[1250] = 3'b010; // x=10, y=31
        pixel_data[1251] = 3'b010; // x=11, y=31
        pixel_data[1252] = 3'b010; // x=12, y=31
        pixel_data[1253] = 3'b010; // x=13, y=31
        pixel_data[1254] = 3'b010; // x=14, y=31
        pixel_data[1255] = 3'b010; // x=15, y=31
        pixel_data[1256] = 3'b010; // x=16, y=31
        pixel_data[1257] = 3'b010; // x=17, y=31
        pixel_data[1258] = 3'b010; // x=18, y=31
        pixel_data[1259] = 3'b010; // x=19, y=31
        pixel_data[1260] = 3'b011; // x=20, y=31
        pixel_data[1261] = 3'b010; // x=21, y=31
        pixel_data[1262] = 3'b011; // x=22, y=31
        pixel_data[1263] = 3'b010; // x=23, y=31
        pixel_data[1264] = 3'b010; // x=24, y=31
        pixel_data[1265] = 3'b010; // x=25, y=31
        pixel_data[1266] = 3'b010; // x=26, y=31
        pixel_data[1267] = 3'b010; // x=27, y=31
        pixel_data[1268] = 3'b010; // x=28, y=31
        pixel_data[1269] = 3'b010; // x=29, y=31
        pixel_data[1270] = 3'b010; // x=30, y=31
        pixel_data[1271] = 3'b011; // x=31, y=31
        pixel_data[1272] = 3'b010; // x=32, y=31
        pixel_data[1273] = 3'b010; // x=33, y=31
        pixel_data[1274] = 3'b010; // x=34, y=31
        pixel_data[1275] = 3'b010; // x=35, y=31
        pixel_data[1276] = 3'b010; // x=36, y=31
        pixel_data[1277] = 3'b010; // x=37, y=31
        pixel_data[1278] = 3'b010; // x=38, y=31
        pixel_data[1279] = 3'b010; // x=39, y=31
        pixel_data[1280] = 3'b010; // x=0, y=32
        pixel_data[1281] = 3'b010; // x=1, y=32
        pixel_data[1282] = 3'b010; // x=2, y=32
        pixel_data[1283] = 3'b010; // x=3, y=32
        pixel_data[1284] = 3'b010; // x=4, y=32
        pixel_data[1285] = 3'b010; // x=5, y=32
        pixel_data[1286] = 3'b010; // x=6, y=32
        pixel_data[1287] = 3'b010; // x=7, y=32
        pixel_data[1288] = 3'b010; // x=8, y=32
        pixel_data[1289] = 3'b010; // x=9, y=32
        pixel_data[1290] = 3'b010; // x=10, y=32
        pixel_data[1291] = 3'b010; // x=11, y=32
        pixel_data[1292] = 3'b010; // x=12, y=32
        pixel_data[1293] = 3'b010; // x=13, y=32
        pixel_data[1294] = 3'b010; // x=14, y=32
        pixel_data[1295] = 3'b010; // x=15, y=32
        pixel_data[1296] = 3'b010; // x=16, y=32
        pixel_data[1297] = 3'b010; // x=17, y=32
        pixel_data[1298] = 3'b010; // x=18, y=32
        pixel_data[1299] = 3'b010; // x=19, y=32
        pixel_data[1300] = 3'b010; // x=20, y=32
        pixel_data[1301] = 3'b011; // x=21, y=32
        pixel_data[1302] = 3'b010; // x=22, y=32
        pixel_data[1303] = 3'b010; // x=23, y=32
        pixel_data[1304] = 3'b010; // x=24, y=32
        pixel_data[1305] = 3'b010; // x=25, y=32
        pixel_data[1306] = 3'b010; // x=26, y=32
        pixel_data[1307] = 3'b010; // x=27, y=32
        pixel_data[1308] = 3'b010; // x=28, y=32
        pixel_data[1309] = 3'b010; // x=29, y=32
        pixel_data[1310] = 3'b010; // x=30, y=32
        pixel_data[1311] = 3'b010; // x=31, y=32
        pixel_data[1312] = 3'b011; // x=32, y=32
        pixel_data[1313] = 3'b010; // x=33, y=32
        pixel_data[1314] = 3'b010; // x=34, y=32
        pixel_data[1315] = 3'b010; // x=35, y=32
        pixel_data[1316] = 3'b010; // x=36, y=32
        pixel_data[1317] = 3'b010; // x=37, y=32
        pixel_data[1318] = 3'b010; // x=38, y=32
        pixel_data[1319] = 3'b010; // x=39, y=32
        pixel_data[1320] = 3'b010; // x=0, y=33
        pixel_data[1321] = 3'b011; // x=1, y=33
        pixel_data[1322] = 3'b010; // x=2, y=33
        pixel_data[1323] = 3'b010; // x=3, y=33
        pixel_data[1324] = 3'b010; // x=4, y=33
        pixel_data[1325] = 3'b010; // x=5, y=33
        pixel_data[1326] = 3'b010; // x=6, y=33
        pixel_data[1327] = 3'b010; // x=7, y=33
        pixel_data[1328] = 3'b010; // x=8, y=33
        pixel_data[1329] = 3'b010; // x=9, y=33
        pixel_data[1330] = 3'b010; // x=10, y=33
        pixel_data[1331] = 3'b011; // x=11, y=33
        pixel_data[1332] = 3'b010; // x=12, y=33
        pixel_data[1333] = 3'b010; // x=13, y=33
        pixel_data[1334] = 3'b010; // x=14, y=33
        pixel_data[1335] = 3'b010; // x=15, y=33
        pixel_data[1336] = 3'b010; // x=16, y=33
        pixel_data[1337] = 3'b010; // x=17, y=33
        pixel_data[1338] = 3'b010; // x=18, y=33
        pixel_data[1339] = 3'b010; // x=19, y=33
        pixel_data[1340] = 3'b010; // x=20, y=33
        pixel_data[1341] = 3'b010; // x=21, y=33
        pixel_data[1342] = 3'b011; // x=22, y=33
        pixel_data[1343] = 3'b010; // x=23, y=33
        pixel_data[1344] = 3'b010; // x=24, y=33
        pixel_data[1345] = 3'b010; // x=25, y=33
        pixel_data[1346] = 3'b010; // x=26, y=33
        pixel_data[1347] = 3'b010; // x=27, y=33
        pixel_data[1348] = 3'b010; // x=28, y=33
        pixel_data[1349] = 3'b010; // x=29, y=33
        pixel_data[1350] = 3'b010; // x=30, y=33
        pixel_data[1351] = 3'b011; // x=31, y=33
        pixel_data[1352] = 3'b010; // x=32, y=33
        pixel_data[1353] = 3'b011; // x=33, y=33
        pixel_data[1354] = 3'b010; // x=34, y=33
        pixel_data[1355] = 3'b010; // x=35, y=33
        pixel_data[1356] = 3'b010; // x=36, y=33
        pixel_data[1357] = 3'b010; // x=37, y=33
        pixel_data[1358] = 3'b010; // x=38, y=33
        pixel_data[1359] = 3'b010; // x=39, y=33
        pixel_data[1360] = 3'b010; // x=0, y=34
        pixel_data[1361] = 3'b010; // x=1, y=34
        pixel_data[1362] = 3'b010; // x=2, y=34
        pixel_data[1363] = 3'b010; // x=3, y=34
        pixel_data[1364] = 3'b010; // x=4, y=34
        pixel_data[1365] = 3'b010; // x=5, y=34
        pixel_data[1366] = 3'b010; // x=6, y=34
        pixel_data[1367] = 3'b010; // x=7, y=34
        pixel_data[1368] = 3'b011; // x=8, y=34
        pixel_data[1369] = 3'b011; // x=9, y=34
        pixel_data[1370] = 3'b010; // x=10, y=34
        pixel_data[1371] = 3'b010; // x=11, y=34
        pixel_data[1372] = 3'b011; // x=12, y=34
        pixel_data[1373] = 3'b010; // x=13, y=34
        pixel_data[1374] = 3'b010; // x=14, y=34
        pixel_data[1375] = 3'b010; // x=15, y=34
        pixel_data[1376] = 3'b010; // x=16, y=34
        pixel_data[1377] = 3'b010; // x=17, y=34
        pixel_data[1378] = 3'b010; // x=18, y=34
        pixel_data[1379] = 3'b010; // x=19, y=34
        pixel_data[1380] = 3'b010; // x=20, y=34
        pixel_data[1381] = 3'b010; // x=21, y=34
        pixel_data[1382] = 3'b010; // x=22, y=34
        pixel_data[1383] = 3'b011; // x=23, y=34
        pixel_data[1384] = 3'b010; // x=24, y=34
        pixel_data[1385] = 3'b010; // x=25, y=34
        pixel_data[1386] = 3'b010; // x=26, y=34
        pixel_data[1387] = 3'b010; // x=27, y=34
        pixel_data[1388] = 3'b010; // x=28, y=34
        pixel_data[1389] = 3'b010; // x=29, y=34
        pixel_data[1390] = 3'b011; // x=30, y=34
        pixel_data[1391] = 3'b010; // x=31, y=34
        pixel_data[1392] = 3'b010; // x=32, y=34
        pixel_data[1393] = 3'b010; // x=33, y=34
        pixel_data[1394] = 3'b011; // x=34, y=34
        pixel_data[1395] = 3'b010; // x=35, y=34
        pixel_data[1396] = 3'b010; // x=36, y=34
        pixel_data[1397] = 3'b010; // x=37, y=34
        pixel_data[1398] = 3'b010; // x=38, y=34
        pixel_data[1399] = 3'b010; // x=39, y=34
        pixel_data[1400] = 3'b010; // x=0, y=35
        pixel_data[1401] = 3'b010; // x=1, y=35
        pixel_data[1402] = 3'b010; // x=2, y=35
        pixel_data[1403] = 3'b010; // x=3, y=35
        pixel_data[1404] = 3'b010; // x=4, y=35
        pixel_data[1405] = 3'b010; // x=5, y=35
        pixel_data[1406] = 3'b010; // x=6, y=35
        pixel_data[1407] = 3'b010; // x=7, y=35
        pixel_data[1408] = 3'b010; // x=8, y=35
        pixel_data[1409] = 3'b010; // x=9, y=35
        pixel_data[1410] = 3'b010; // x=10, y=35
        pixel_data[1411] = 3'b010; // x=11, y=35
        pixel_data[1412] = 3'b010; // x=12, y=35
        pixel_data[1413] = 3'b011; // x=13, y=35
        pixel_data[1414] = 3'b010; // x=14, y=35
        pixel_data[1415] = 3'b010; // x=15, y=35
        pixel_data[1416] = 3'b010; // x=16, y=35
        pixel_data[1417] = 3'b010; // x=17, y=35
        pixel_data[1418] = 3'b011; // x=18, y=35
        pixel_data[1419] = 3'b010; // x=19, y=35
        pixel_data[1420] = 3'b010; // x=20, y=35
        pixel_data[1421] = 3'b010; // x=21, y=35
        pixel_data[1422] = 3'b010; // x=22, y=35
        pixel_data[1423] = 3'b010; // x=23, y=35
        pixel_data[1424] = 3'b011; // x=24, y=35
        pixel_data[1425] = 3'b010; // x=25, y=35
        pixel_data[1426] = 3'b010; // x=26, y=35
        pixel_data[1427] = 3'b010; // x=27, y=35
        pixel_data[1428] = 3'b010; // x=28, y=35
        pixel_data[1429] = 3'b011; // x=29, y=35
        pixel_data[1430] = 3'b010; // x=30, y=35
        pixel_data[1431] = 3'b010; // x=31, y=35
        pixel_data[1432] = 3'b010; // x=32, y=35
        pixel_data[1433] = 3'b010; // x=33, y=35
        pixel_data[1434] = 3'b010; // x=34, y=35
        pixel_data[1435] = 3'b011; // x=35, y=35
        pixel_data[1436] = 3'b010; // x=36, y=35
        pixel_data[1437] = 3'b010; // x=37, y=35
        pixel_data[1438] = 3'b010; // x=38, y=35
        pixel_data[1439] = 3'b010; // x=39, y=35
        pixel_data[1440] = 3'b010; // x=0, y=36
        pixel_data[1441] = 3'b010; // x=1, y=36
        pixel_data[1442] = 3'b010; // x=2, y=36
        pixel_data[1443] = 3'b011; // x=3, y=36
        pixel_data[1444] = 3'b010; // x=4, y=36
        pixel_data[1445] = 3'b011; // x=5, y=36
        pixel_data[1446] = 3'b011; // x=6, y=36
        pixel_data[1447] = 3'b010; // x=7, y=36
        pixel_data[1448] = 3'b010; // x=8, y=36
        pixel_data[1449] = 3'b010; // x=9, y=36
        pixel_data[1450] = 3'b010; // x=10, y=36
        pixel_data[1451] = 3'b010; // x=11, y=36
        pixel_data[1452] = 3'b010; // x=12, y=36
        pixel_data[1453] = 3'b010; // x=13, y=36
        pixel_data[1454] = 3'b011; // x=14, y=36
        pixel_data[1455] = 3'b010; // x=15, y=36
        pixel_data[1456] = 3'b011; // x=16, y=36
        pixel_data[1457] = 3'b010; // x=17, y=36
        pixel_data[1458] = 3'b000; // x=18, y=36
        pixel_data[1459] = 3'b000; // x=19, y=36
        pixel_data[1460] = 3'b000; // x=20, y=36
        pixel_data[1461] = 3'b000; // x=21, y=36
        pixel_data[1462] = 3'b000; // x=22, y=36
        pixel_data[1463] = 3'b010; // x=23, y=36
        pixel_data[1464] = 3'b010; // x=24, y=36
        pixel_data[1465] = 3'b010; // x=25, y=36
        pixel_data[1466] = 3'b010; // x=26, y=36
        pixel_data[1467] = 3'b011; // x=27, y=36
        pixel_data[1468] = 3'b011; // x=28, y=36
        pixel_data[1469] = 3'b010; // x=29, y=36
        pixel_data[1470] = 3'b010; // x=30, y=36
        pixel_data[1471] = 3'b010; // x=31, y=36
        pixel_data[1472] = 3'b010; // x=32, y=36
        pixel_data[1473] = 3'b010; // x=33, y=36
        pixel_data[1474] = 3'b010; // x=34, y=36
        pixel_data[1475] = 3'b010; // x=35, y=36
        pixel_data[1476] = 3'b010; // x=36, y=36
        pixel_data[1477] = 3'b010; // x=37, y=36
        pixel_data[1478] = 3'b011; // x=38, y=36
        pixel_data[1479] = 3'b011; // x=39, y=36
        pixel_data[1480] = 3'b010; // x=0, y=37
        pixel_data[1481] = 3'b010; // x=1, y=37
        pixel_data[1482] = 3'b010; // x=2, y=37
        pixel_data[1483] = 3'b010; // x=3, y=37
        pixel_data[1484] = 3'b011; // x=4, y=37
        pixel_data[1485] = 3'b011; // x=5, y=37
        pixel_data[1486] = 3'b011; // x=6, y=37
        pixel_data[1487] = 3'b010; // x=7, y=37
        pixel_data[1488] = 3'b010; // x=8, y=37
        pixel_data[1489] = 3'b010; // x=9, y=37
        pixel_data[1490] = 3'b010; // x=10, y=37
        pixel_data[1491] = 3'b010; // x=11, y=37
        pixel_data[1492] = 3'b010; // x=12, y=37
        pixel_data[1493] = 3'b010; // x=13, y=37
        pixel_data[1494] = 3'b010; // x=14, y=37
        pixel_data[1495] = 3'b011; // x=15, y=37
        pixel_data[1496] = 3'b011; // x=16, y=37
        pixel_data[1497] = 3'b100; // x=17, y=37
        pixel_data[1498] = 3'b101; // x=18, y=37
        pixel_data[1499] = 3'b101; // x=19, y=37
        pixel_data[1500] = 3'b101; // x=20, y=37
        pixel_data[1501] = 3'b101; // x=21, y=37
        pixel_data[1502] = 3'b100; // x=22, y=37
        pixel_data[1503] = 3'b011; // x=23, y=37
        pixel_data[1504] = 3'b010; // x=24, y=37
        pixel_data[1505] = 3'b010; // x=25, y=37
        pixel_data[1506] = 3'b011; // x=26, y=37
        pixel_data[1507] = 3'b011; // x=27, y=37
        pixel_data[1508] = 3'b011; // x=28, y=37
        pixel_data[1509] = 3'b010; // x=29, y=37
        pixel_data[1510] = 3'b010; // x=30, y=37
        pixel_data[1511] = 3'b010; // x=31, y=37
        pixel_data[1512] = 3'b010; // x=32, y=37
        pixel_data[1513] = 3'b010; // x=33, y=37
        pixel_data[1514] = 3'b010; // x=34, y=37
        pixel_data[1515] = 3'b010; // x=35, y=37
        pixel_data[1516] = 3'b010; // x=36, y=37
        pixel_data[1517] = 3'b011; // x=37, y=37
        pixel_data[1518] = 3'b011; // x=38, y=37
        pixel_data[1519] = 3'b011; // x=39, y=37
        pixel_data[1520] = 3'b010; // x=0, y=38
        pixel_data[1521] = 3'b010; // x=1, y=38
        pixel_data[1522] = 3'b010; // x=2, y=38
        pixel_data[1523] = 3'b011; // x=3, y=38
        pixel_data[1524] = 3'b011; // x=4, y=38
        pixel_data[1525] = 3'b011; // x=5, y=38
        pixel_data[1526] = 3'b011; // x=6, y=38
        pixel_data[1527] = 3'b010; // x=7, y=38
        pixel_data[1528] = 3'b010; // x=8, y=38
        pixel_data[1529] = 3'b010; // x=9, y=38
        pixel_data[1530] = 3'b010; // x=10, y=38
        pixel_data[1531] = 3'b010; // x=11, y=38
        pixel_data[1532] = 3'b010; // x=12, y=38
        pixel_data[1533] = 3'b010; // x=13, y=38
        pixel_data[1534] = 3'b011; // x=14, y=38
        pixel_data[1535] = 3'b011; // x=15, y=38
        pixel_data[1536] = 3'b011; // x=16, y=38
        pixel_data[1537] = 3'b101; // x=17, y=38
        pixel_data[1538] = 3'b101; // x=18, y=38
        pixel_data[1539] = 3'b101; // x=19, y=38
        pixel_data[1540] = 3'b101; // x=20, y=38
        pixel_data[1541] = 3'b101; // x=21, y=38
        pixel_data[1542] = 3'b100; // x=22, y=38
        pixel_data[1543] = 3'b011; // x=23, y=38
        pixel_data[1544] = 3'b001; // x=24, y=38
        pixel_data[1545] = 3'b011; // x=25, y=38
        pixel_data[1546] = 3'b011; // x=26, y=38
        pixel_data[1547] = 3'b011; // x=27, y=38
        pixel_data[1548] = 3'b010; // x=28, y=38
        pixel_data[1549] = 3'b010; // x=29, y=38
        pixel_data[1550] = 3'b010; // x=30, y=38
        pixel_data[1551] = 3'b010; // x=31, y=38
        pixel_data[1552] = 3'b010; // x=32, y=38
        pixel_data[1553] = 3'b010; // x=33, y=38
        pixel_data[1554] = 3'b010; // x=34, y=38
        pixel_data[1555] = 3'b010; // x=35, y=38
        pixel_data[1556] = 3'b011; // x=36, y=38
        pixel_data[1557] = 3'b011; // x=37, y=38
        pixel_data[1558] = 3'b011; // x=38, y=38
        pixel_data[1559] = 3'b010; // x=39, y=38
        pixel_data[1560] = 3'b010; // x=0, y=39
        pixel_data[1561] = 3'b010; // x=1, y=39
        pixel_data[1562] = 3'b010; // x=2, y=39
        pixel_data[1563] = 3'b011; // x=3, y=39
        pixel_data[1564] = 3'b011; // x=4, y=39
        pixel_data[1565] = 3'b010; // x=5, y=39
        pixel_data[1566] = 3'b011; // x=6, y=39
        pixel_data[1567] = 3'b010; // x=7, y=39
        pixel_data[1568] = 3'b010; // x=8, y=39
        pixel_data[1569] = 3'b010; // x=9, y=39
        pixel_data[1570] = 3'b010; // x=10, y=39
        pixel_data[1571] = 3'b010; // x=11, y=39
        pixel_data[1572] = 3'b010; // x=12, y=39
        pixel_data[1573] = 3'b010; // x=13, y=39
        pixel_data[1574] = 3'b011; // x=14, y=39
        pixel_data[1575] = 3'b011; // x=15, y=39
        pixel_data[1576] = 3'b010; // x=16, y=39
        pixel_data[1577] = 3'b000; // x=17, y=39
        pixel_data[1578] = 3'b000; // x=18, y=39
        pixel_data[1579] = 3'b000; // x=19, y=39
        pixel_data[1580] = 3'b000; // x=20, y=39
        pixel_data[1581] = 3'b000; // x=21, y=39
        pixel_data[1582] = 3'b000; // x=22, y=39
        pixel_data[1583] = 3'b010; // x=23, y=39
        pixel_data[1584] = 3'b010; // x=24, y=39
        pixel_data[1585] = 3'b011; // x=25, y=39
        pixel_data[1586] = 3'b011; // x=26, y=39
        pixel_data[1587] = 3'b011; // x=27, y=39
        pixel_data[1588] = 3'b010; // x=28, y=39
        pixel_data[1589] = 3'b010; // x=29, y=39
        pixel_data[1590] = 3'b010; // x=30, y=39
        pixel_data[1591] = 3'b010; // x=31, y=39
        pixel_data[1592] = 3'b010; // x=32, y=39
        pixel_data[1593] = 3'b010; // x=33, y=39
        pixel_data[1594] = 3'b010; // x=34, y=39
        pixel_data[1595] = 3'b011; // x=35, y=39
        pixel_data[1596] = 3'b011; // x=36, y=39
        pixel_data[1597] = 3'b011; // x=37, y=39
        pixel_data[1598] = 3'b010; // x=38, y=39
        pixel_data[1599] = 3'b011; // x=39, y=39
    end
endmodule
